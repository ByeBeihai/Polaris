module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [8:0]  io_rreq_bits_setIdx,
  output [27:0] io_rresp_data_0_tag,
  output [1:0]  io_rresp_data_0__type,
  output [38:0] io_rresp_data_0_target,
  output [2:0]  io_rresp_data_0_brIdx,
  output        io_rresp_data_0_valid,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [27:0] io_wreq_bits_data_tag,
  input  [1:0]  io_wreq_bits_data__type,
  input  [38:0] io_wreq_bits_data_target,
  input  [2:0]  io_wreq_bits_data_brIdx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  reg  REG; // @[SRAMTemplate.scala 80:30]
  reg [8:0] value; // @[Counter.scala 60:40]
  wire  wrap_wrap = value == 9'h1ff; // @[Counter.scala 72:24]
  wire [8:0] _wrap_value_T_1 = value + 9'h1; // @[Counter.scala 76:24]
  wire  wrap = REG & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = wrap ? 1'h0 : REG; // @[SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  wire  _T = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = REG ? value : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [72:0] _T_1 = {io_wreq_bits_data_tag,io_wreq_bits_data__type,io_wreq_bits_data_target,io_wreq_bits_data_brIdx
    ,1'h1}; // @[SRAMTemplate.scala 92:78]
  reg  REG_1; // @[Hold.scala 28:106]
  reg [72:0] r_0; // @[Reg.scala 27:20]
  wire [72:0] _GEN_14 = REG_1 ? array_RW0_rdata_0 : r_0; // @[Reg.scala 28:19 27:20 28:23]
  array array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_rdata_0(array_RW0_rdata_0)
  );
  assign io_rreq_ready = ~REG & _T; // @[SRAMTemplate.scala 101:33]
  assign io_rresp_data_0_tag = _GEN_14[72:45]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0__type = _GEN_14[44:43]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_target = _GEN_14[42:4]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_brIdx = _GEN_14[3:1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_valid = _GEN_14[0]; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = REG ? 73'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_en = realRen | wen;
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[Counter.scala 60:40]
      value <= 9'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      value <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    REG_1 <= io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
    if (reset) begin // @[Reg.scala 27:20]
      r_0 <= 73'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_0 <= array_RW0_rdata_0; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {3{`RANDOM}};
  r_0 = _RAND_3[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid,
  input  [38:0] io_in_pc_bits,
  output [38:0] io_out_target,
  output        io_out_valid,
  input         io_flush,
  output [2:0]  io_brIdx,
  output        io_crosslineJump,
  input         MOUFlushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[BPU.scala 335:19]
  wire  btb_reset; // @[BPU.scala 335:19]
  wire  btb_io_rreq_ready; // @[BPU.scala 335:19]
  wire  btb_io_rreq_valid; // @[BPU.scala 335:19]
  wire [8:0] btb_io_rreq_bits_setIdx; // @[BPU.scala 335:19]
  wire [27:0] btb_io_rresp_data_0_tag; // @[BPU.scala 335:19]
  wire [1:0] btb_io_rresp_data_0__type; // @[BPU.scala 335:19]
  wire [38:0] btb_io_rresp_data_0_target; // @[BPU.scala 335:19]
  wire [2:0] btb_io_rresp_data_0_brIdx; // @[BPU.scala 335:19]
  wire  btb_io_rresp_data_0_valid; // @[BPU.scala 335:19]
  wire  btb_io_wreq_valid; // @[BPU.scala 335:19]
  wire [8:0] btb_io_wreq_bits_setIdx; // @[BPU.scala 335:19]
  wire [27:0] btb_io_wreq_bits_data_tag; // @[BPU.scala 335:19]
  wire [1:0] btb_io_wreq_bits_data__type; // @[BPU.scala 335:19]
  wire [38:0] btb_io_wreq_bits_data_target; // @[BPU.scala 335:19]
  wire [2:0] btb_io_wreq_bits_data_brIdx; // @[BPU.scala 335:19]
  reg [1:0] pht [0:511]; // @[BPU.scala 369:16]
  wire  pht_MPORT_en; // @[BPU.scala 369:16]
  wire [8:0] pht_MPORT_addr; // @[BPU.scala 369:16]
  wire [1:0] pht_MPORT_data; // @[BPU.scala 369:16]
  wire  pht_MPORT_2_en; // @[BPU.scala 369:16]
  wire [8:0] pht_MPORT_2_addr; // @[BPU.scala 369:16]
  wire [1:0] pht_MPORT_2_data; // @[BPU.scala 369:16]
  wire  pht_MPORT_5_en; // @[BPU.scala 369:16]
  wire [8:0] pht_MPORT_5_addr; // @[BPU.scala 369:16]
  wire [1:0] pht_MPORT_5_data; // @[BPU.scala 369:16]
  wire [1:0] pht_MPORT_3_data; // @[BPU.scala 369:16]
  wire [8:0] pht_MPORT_3_addr; // @[BPU.scala 369:16]
  wire  pht_MPORT_3_mask; // @[BPU.scala 369:16]
  wire  pht_MPORT_3_en; // @[BPU.scala 369:16]
  reg [38:0] ras [0:15]; // @[BPU.scala 375:16]
  wire  ras_MPORT_1_en; // @[BPU.scala 375:16]
  wire [3:0] ras_MPORT_1_addr; // @[BPU.scala 375:16]
  wire [38:0] ras_MPORT_1_data; // @[BPU.scala 375:16]
  wire [38:0] ras_MPORT_4_data; // @[BPU.scala 375:16]
  wire [3:0] ras_MPORT_4_addr; // @[BPU.scala 375:16]
  wire  ras_MPORT_4_mask; // @[BPU.scala 375:16]
  wire  ras_MPORT_4_en; // @[BPU.scala 375:16]
  reg  flush; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = io_flush | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg [38:0] pcLatch; // @[Reg.scala 15:16]
  wire [27:0] btbRead_tag = btb_io_rresp_data_0_tag; // @[BPU.scala 348:21 349:11]
  wire  btbRead_valid = btb_io_rresp_data_0_valid; // @[BPU.scala 348:21 349:11]
  wire  _T_23 = btb_io_rreq_ready & btb_io_rreq_valid; // @[Decoupled.scala 40:37]
  reg  REG_1; // @[BPU.scala 353:93]
  wire [2:0] btbRead_brIdx = btb_io_rresp_data_0_brIdx; // @[BPU.scala 348:21 349:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:11] & ~flush & REG_1 & ~(pcLatch[1] & btbRead_brIdx[0]); // @[BPU.scala 353:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 360:40]
  reg  phtTaken; // @[Reg.scala 15:16]
  reg [3:0] value; // @[Counter.scala 60:40]
  reg [38:0] rasTarget; // @[Reg.scala 15:16]
  wire  _T_40 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[BPU.scala 399:46]
  wire  _T_43 = ~bpuUpdateReq_pc[1]; // @[BPU.scala 399:72]
  wire [1:0] hi = {_T_40,bpuUpdateReq_pc[1]}; // @[Cat.scala 30:58]
  reg [1:0] cnt; // @[BPU.scala 421:20]
  reg  reqLatch_valid; // @[BPU.scala 422:25]
  reg [38:0] reqLatch_pc; // @[BPU.scala 422:25]
  reg  reqLatch_actualTaken; // @[BPU.scala 422:25]
  reg [6:0] reqLatch_fuOpType; // @[BPU.scala 422:25]
  wire  _T_70 = ~reqLatch_fuOpType[3]; // @[ALU.scala 70:30]
  wire  _T_71 = reqLatch_valid & _T_70; // @[BPU.scala 423:24]
  wire [1:0] _T_73 = cnt + 2'h1; // @[BPU.scala 425:33]
  wire [1:0] _T_75 = cnt - 2'h1; // @[BPU.scala 425:44]
  wire  _T_82 = reqLatch_actualTaken & cnt != 2'h3 | ~reqLatch_actualTaken & cnt != 2'h0; // @[BPU.scala 426:44]
  wire  _T_93 = bpuUpdateReq_fuOpType == 7'h5c; // @[BPU.scala 433:24]
  wire [3:0] _T_95 = value + 4'h1; // @[BPU.scala 434:26]
  wire [38:0] _T_97 = bpuUpdateReq_pc + 39'h2; // @[BPU.scala 434:55]
  wire [38:0] _T_99 = bpuUpdateReq_pc + 39'h4; // @[BPU.scala 434:69]
  wire  _T_102 = value == 4'h0; // @[BPU.scala 439:21]
  wire [3:0] _value_T_4 = value - 4'h1; // @[BPU.scala 442:53]
  wire [3:0] _value_T_5 = _T_102 ? 4'h0 : _value_T_4; // @[BPU.scala 442:22]
  wire [1:0] btbRead__type = btb_io_rresp_data_0__type; // @[BPU.scala 348:21 349:11]
  wire [38:0] btbRead_target = btb_io_rresp_data_0_target; // @[BPU.scala 348:21 349:11]
  wire [1:0] _T_106 = io_out_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_107 = {1'h1,crosslineJump,_T_106}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_28 = {{1'd0}, btbRead_brIdx}; // @[BPU.scala 449:30]
  wire [3:0] _T_108 = _GEN_28 & _T_107; // @[BPU.scala 449:30]
  wire  _T_112 = btbRead__type == 2'h0 ? phtTaken : rasTarget != 39'h0; // @[BPU.scala 450:32]
  SRAMTemplate btb ( // @[BPU.scala 335:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_rreq_ready(btb_io_rreq_ready),
    .io_rreq_valid(btb_io_rreq_valid),
    .io_rreq_bits_setIdx(btb_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(btb_io_rresp_data_0_tag),
    .io_rresp_data_0__type(btb_io_rresp_data_0__type),
    .io_rresp_data_0_target(btb_io_rresp_data_0_target),
    .io_rresp_data_0_brIdx(btb_io_rresp_data_0_brIdx),
    .io_rresp_data_0_valid(btb_io_rresp_data_0_valid),
    .io_wreq_valid(btb_io_wreq_valid),
    .io_wreq_bits_setIdx(btb_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(btb_io_wreq_bits_data_tag),
    .io_wreq_bits_data__type(btb_io_wreq_bits_data__type),
    .io_wreq_bits_data_target(btb_io_wreq_bits_data_target),
    .io_wreq_bits_data_brIdx(btb_io_wreq_bits_data_brIdx)
  );
  assign pht_MPORT_en = 1'h1;
  assign pht_MPORT_addr = io_in_pc_bits[10:2];
  assign pht_MPORT_data = pht[pht_MPORT_addr]; // @[BPU.scala 369:16]
  assign pht_MPORT_2_en = 1'h1;
  assign pht_MPORT_2_addr = bpuUpdateReq_pc[10:2];
  assign pht_MPORT_2_data = pht[pht_MPORT_2_addr]; // @[BPU.scala 369:16]
  assign pht_MPORT_5_en = 1'h1;
  assign pht_MPORT_5_addr = io_in_pc_bits[10:2];
  assign pht_MPORT_5_data = pht[pht_MPORT_5_addr]; // @[BPU.scala 369:16]
  assign pht_MPORT_3_data = reqLatch_actualTaken ? _T_73 : _T_75;
  assign pht_MPORT_3_addr = reqLatch_pc[10:2];
  assign pht_MPORT_3_mask = 1'h1;
  assign pht_MPORT_3_en = _T_71 & _T_82;
  assign ras_MPORT_1_en = 1'h1;
  assign ras_MPORT_1_addr = value;
  assign ras_MPORT_1_data = ras[ras_MPORT_1_addr]; // @[BPU.scala 375:16]
  assign ras_MPORT_4_data = bpuUpdateReq_isRVC ? _T_97 : _T_99;
  assign ras_MPORT_4_addr = value + 4'h1;
  assign ras_MPORT_4_mask = 1'h1;
  assign ras_MPORT_4_en = bpuUpdateReq_valid & _T_93;
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[BPU.scala 446:23]
  assign io_out_valid = btbHit & _T_112; // @[BPU.scala 450:26]
  assign io_brIdx = _T_108[2:0]; // @[BPU.scala 449:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 360:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[BPU.scala 341:29]
  assign btb_io_rreq_valid = io_in_pc_valid; // @[BPU.scala 344:22]
  assign btb_io_rreq_bits_setIdx = io_in_pc_bits[10:2]; // @[BPU.scala 35:65]
  assign btb_io_wreq_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[BPU.scala 407:43]
  assign btb_io_wreq_bits_setIdx = bpuUpdateReq_pc[10:2]; // @[BPU.scala 35:65]
  assign btb_io_wreq_bits_data_tag = bpuUpdateReq_pc[38:11]; // @[BPU.scala 35:65]
  assign btb_io_wreq_bits_data__type = bpuUpdateReq_btbType; // @[BPU.scala 409:26]
  assign btb_io_wreq_bits_data_target = bpuUpdateReq_actualTarget; // @[BPU.scala 409:26]
  assign btb_io_wreq_bits_data_brIdx = {hi,_T_43}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (pht_MPORT_3_en & pht_MPORT_3_mask) begin
      pht[pht_MPORT_3_addr] <= pht_MPORT_3_data; // @[BPU.scala 369:16]
    end
    if (ras_MPORT_4_en & ras_MPORT_4_mask) begin
      ras[ras_MPORT_4_addr] <= ras_MPORT_4_data; // @[BPU.scala 375:16]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      flush <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (io_in_pc_valid) begin // @[Reg.scala 16:19]
      pcLatch <= io_in_pc_bits; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[BPU.scala 353:93]
      REG_1 <= 1'h0; // @[BPU.scala 353:93]
    end else begin
      REG_1 <= _T_23; // @[BPU.scala 353:93]
    end
    if (io_in_pc_valid) begin // @[Reg.scala 16:19]
      phtTaken <= pht_MPORT_data[1]; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 4'h0; // @[Counter.scala 60:40]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 432:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 433:45]
        value <= _T_95; // @[BPU.scala 436:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[BPU.scala 438:48]
        value <= _value_T_5; // @[BPU.scala 442:16]
      end
    end
    if (io_in_pc_valid) begin // @[Reg.scala 16:19]
      rasTarget <= ras_MPORT_1_data; // @[Reg.scala 16:23]
    end
    cnt <= pht_MPORT_2_data; // @[BPU.scala 421:20]
    reqLatch_valid <= bpuUpdateReq_valid; // @[BPU.scala 422:25]
    reqLatch_pc <= bpuUpdateReq_pc; // @[BPU.scala 422:25]
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken; // @[BPU.scala 422:25]
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType; // @[BPU.scala 422:25]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    pht[initvar] = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_1[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  flush = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  pcLatch = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  phtTaken = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[3:0];
  _RAND_7 = {2{`RANDOM}};
  rasTarget = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  cnt = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reqLatch_valid = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  reqLatch_pc = _RAND_10[38:0];
  _RAND_11 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_12[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [81:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [81:0] io_imem_resp_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input         flushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[IFU.scala 107:19]
  wire  bp1_reset; // @[IFU.scala 107:19]
  wire  bp1_io_in_pc_valid; // @[IFU.scala 107:19]
  wire [38:0] bp1_io_in_pc_bits; // @[IFU.scala 107:19]
  wire [38:0] bp1_io_out_target; // @[IFU.scala 107:19]
  wire  bp1_io_out_valid; // @[IFU.scala 107:19]
  wire  bp1_io_flush; // @[IFU.scala 107:19]
  wire [2:0] bp1_io_brIdx; // @[IFU.scala 107:19]
  wire  bp1_io_crosslineJump; // @[IFU.scala 107:19]
  wire  bp1_MOUFlushICache; // @[IFU.scala 107:19]
  wire  bp1_bpuUpdateReq_valid; // @[IFU.scala 107:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[IFU.scala 107:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[IFU.scala 107:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[IFU.scala 107:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[IFU.scala 107:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[IFU.scala 107:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[IFU.scala 107:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[IFU.scala 107:19]
  wire  bp1_MOUFlushTLB; // @[IFU.scala 107:19]
  reg [38:0] pc; // @[IFU.scala 103:19]
  wire  _T = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire  pcUpdate = io_redirect_valid | _T; // @[IFU.scala 104:36]
  wire [38:0] _T_3 = pc + 39'h2; // @[IFU.scala 105:28]
  wire [38:0] _T_5 = pc + 39'h4; // @[IFU.scala 105:38]
  wire [38:0] snpc = pc[1] ? _T_3 : _T_5; // @[IFU.scala 105:17]
  reg  crosslineJumpLatch; // @[IFU.scala 110:35]
  reg [38:0] crosslineJumpTarget; // @[Reg.scala 15:16]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[IFU.scala 119:17]
  wire [38:0] _T_11 = bp1_io_out_valid ? pnpc : snpc; // @[IFU.scala 122:104]
  wire [38:0] _T_12 = crosslineJumpLatch ? crosslineJumpTarget : _T_11; // @[IFU.scala 122:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 122:16]
  wire  _T_13 = bp1_io_out_valid ? 1'h0 : 1'h1; // @[IFU.scala 123:114]
  wire  _T_15 = crosslineJumpLatch ? 1'h0 : bp1_io_crosslineJump | _T_13; // @[IFU.scala 123:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _T_15; // @[IFU.scala 123:21]
  wire [2:0] _T_16 = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[IFU.scala 131:29]
  wire [42:0] hi = {npcIsSeq,_T_16,npc}; // @[Cat.scala 30:58]
  wire  _T_41 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | REG_1; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_42 = |io_flushVec; // @[IFU.scala 178:37]
  BPU_inorder bp1 ( // @[IFU.scala 107:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .MOUFlushICache(bp1_MOUFlushICache),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[IFU.scala 156:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[Cat.scala 30:58]
  assign io_imem_req_bits_user = {hi,pc}; // @[Cat.scala 30:58]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[IFU.scala 158:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[IFU.scala 175:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[IFU.scala 168:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[IFU.scala 170:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[IFU.scala 171:26]
  assign io_out_bits_exceptionVec_12 = io_ipf; // @[IFU.scala 174:44]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[IFU.scala 172:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[IFU.scala 151:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 122:16]
  assign bp1_io_flush = io_redirect_valid; // @[IFU.scala 140:16]
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_bpuUpdateReq_valid = bpuUpdateReq_valid;
  assign bp1_bpuUpdateReq_pc = bpuUpdateReq_pc;
  assign bp1_bpuUpdateReq_isMissPredict = bpuUpdateReq_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = bpuUpdateReq_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = bpuUpdateReq_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = bpuUpdateReq_fuOpType;
  assign bp1_bpuUpdateReq_btbType = bpuUpdateReq_btbType;
  assign bp1_bpuUpdateReq_isRVC = bpuUpdateReq_isRVC;
  assign bp1_MOUFlushTLB = flushTLB;
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 103:19]
      pc <= 39'h80000000; // @[IFU.scala 103:19]
    end else if (pcUpdate) begin // @[IFU.scala 142:19]
      if (io_redirect_valid) begin // @[IFU.scala 122:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[IFU.scala 122:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= _T_11;
      end
    end
    if (reset) begin // @[IFU.scala 110:35]
      crosslineJumpLatch <= 1'h0; // @[IFU.scala 110:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[IFU.scala 111:34]
      if (bp1_io_flush) begin // @[IFU.scala 112:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (bp1_io_crosslineJump) begin // @[Reg.scala 16:19]
      crosslineJumpTarget <= bp1_io_out_target; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_41) begin // @[StopWatch.scala 31:19]
      REG_1 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_1 <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  output        io_out_bits_crossPageIPFFix,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[NaiveIBF.scala 39:22]
  wire  _T_81 = state == 2'h2; // @[NaiveIBF.scala 90:23]
  wire  _T_82 = state == 2'h3; // @[NaiveIBF.scala 90:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[Cat.scala 30:58]
  reg [15:0] specialInstR; // @[NaiveIBF.scala 66:25]
  wire [31:0] _T_85 = {instIn[15:0],specialInstR}; // @[Cat.scala 30:58]
  wire  _T_1 = state == 2'h0; // @[NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[NaiveIBF.scala 41:21]
  wire  _T_90 = 3'h0 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_94 = _T_90 ? instIn[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_91 = 3'h2 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_95 = _T_91 ? instIn[47:16] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_98 = _T_94 | _T_95; // @[Mux.scala 27:72]
  wire  _T_92 = 3'h4 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_96 = _T_92 ? instIn[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_99 = _T_98 | _T_96; // @[Mux.scala 27:72]
  wire  _T_93 = 3'h6 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_97 = _T_93 ? instIn[79:48] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_100 = _T_99 | _T_97; // @[Mux.scala 27:72]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _T_85 : _T_100; // @[NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[NaiveIBF.scala 34:26]
  wire  _T_3 = pcOffset == 3'h0; // @[NaiveIBF.scala 48:28]
  wire  _T_4 = ~isRVC; // @[NaiveIBF.scala 48:40]
  wire  _T_8 = pcOffset == 3'h4; // @[NaiveIBF.scala 48:72]
  wire  _T_14 = pcOffset == 3'h2; // @[NaiveIBF.scala 48:116]
  wire  _T_19 = pcOffset == 3'h6; // @[NaiveIBF.scala 48:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[NaiveIBF.scala 48:147]
  wire  _T_34 = _T_14 & _T_4; // @[NaiveIBF.scala 51:122]
  wire  _T_36 = ~io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:135]
  wire  rvcNext = _T_3 & (isRVC & ~io_in_bits_brIdx[0]) | _T_8 & (isRVC & ~io_in_bits_brIdx[0]) | _T_14 & _T_4 & ~
    io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:102]
  wire  _T_40 = _T_19 & _T_4; // @[NaiveIBF.scala 52:37]
  wire  rvcSpecial = _T_19 & _T_4 & ~io_in_bits_brIdx[2]; // @[NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _T_40 & io_in_bits_brIdx[2]; // @[NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[NaiveIBF.scala 54:24]
  wire  _T_49 = _T_1 | state == 2'h1; // @[NaiveIBF.scala 57:36]
  wire  flushIFU = (_T_1 | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[NaiveIBF.scala 57:87]
  wire  loadNextInstline = _T_49 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[NaiveIBF.scala 64:23]
  reg [38:0] specialNPCR; // @[NaiveIBF.scala 65:24]
  reg  specialIPFR; // @[NaiveIBF.scala 67:28]
  wire  rvcForceLoadNext = _T_34 & io_in_bits_pnpc[2:0] == 3'h4 & _T_36; // @[NaiveIBF.scala 69:86]
  wire  _T_104 = rvcFinish | rvcNext; // @[NaiveIBF.scala 100:28]
  wire  _T_105 = rvcFinish | rvcForceLoadNext; // @[NaiveIBF.scala 101:28]
  wire [38:0] _T_107 = io_in_bits_pc + 39'h2; // @[NaiveIBF.scala 103:76]
  wire [38:0] _T_109 = io_in_bits_pc + 39'h4; // @[NaiveIBF.scala 103:95]
  wire [38:0] _T_110 = isRVC ? _T_107 : _T_109; // @[NaiveIBF.scala 103:55]
  wire [38:0] _T_111 = rvcFinish ? io_in_bits_pnpc : _T_110; // @[NaiveIBF.scala 103:23]
  wire  _T_112 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_0 = _T_112 & rvcFinish ? 2'h0 : state; // @[NaiveIBF.scala 104:{41,48} 39:22]
  wire [2:0] _T_116 = isRVC ? 3'h2 : 3'h4; // @[NaiveIBF.scala 107:38]
  wire [2:0] _T_118 = pcOffset + _T_116; // @[NaiveIBF.scala 107:33]
  wire [1:0] _GEN_1 = _T_112 & rvcNext ? 2'h1 : _GEN_0; // @[NaiveIBF.scala 105:39 106:17]
  wire [2:0] _GEN_2 = _T_112 & rvcNext ? _T_118 : pcOffsetR; // @[NaiveIBF.scala 105:39 107:21 40:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[NaiveIBF.scala 109:40 110:17]
  wire [38:0] _T_128 = {io_in_bits_pc[38:3],pcOffsetR}; // @[Cat.scala 30:58]
  wire [38:0] _GEN_27 = 2'h3 == state ? specialPCR : 39'h0; // @[NaiveIBF.scala 161:15 98:18]
  wire [38:0] _GEN_32 = 2'h2 == state ? specialPCR : _GEN_27; // @[NaiveIBF.scala 149:15 98:18]
  wire [38:0] _GEN_40 = 2'h1 == state ? _T_128 : _GEN_32; // @[NaiveIBF.scala 126:15 98:18]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[NaiveIBF.scala 102:15 98:18]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[NaiveIBF.scala 109:40 111:22 64:23]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[NaiveIBF.scala 109:40 112:24 66:25]
  wire  _GEN_6 = rvcSpecial & io_in_valid ? io_in_bits_exceptionVec_12 : specialIPFR; // @[NaiveIBF.scala 109:40 113:23 67:28]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[NaiveIBF.scala 115:44 116:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[NaiveIBF.scala 115:44 117:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[NaiveIBF.scala 115:44 118:23 65:24]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[NaiveIBF.scala 115:44 119:24]
  wire  _GEN_11 = rvcSpecialJump & io_in_valid ? io_in_bits_exceptionVec_12 : _GEN_6; // @[NaiveIBF.scala 115:44 120:23]
  wire [38:0] _T_130 = pcOut + 39'h2; // @[NaiveIBF.scala 127:68]
  wire [38:0] _T_132 = pcOut + 39'h4; // @[NaiveIBF.scala 127:79]
  wire [38:0] _T_133 = isRVC ? _T_130 : _T_132; // @[NaiveIBF.scala 127:55]
  wire [38:0] _T_134 = rvcFinish ? io_in_bits_pnpc : _T_133; // @[NaiveIBF.scala 127:23]
  wire [38:0] _T_148 = specialPCR + 39'h4; // @[NaiveIBF.scala 150:31]
  wire [1:0] _GEN_24 = _T_112 ? 2'h1 : state; // @[NaiveIBF.scala 154:28 155:17 39:22]
  wire [2:0] _GEN_25 = _T_112 ? 3'h2 : pcOffsetR; // @[NaiveIBF.scala 154:28 156:21 40:26]
  wire [1:0] _GEN_26 = _T_112 ? 2'h0 : state; // @[NaiveIBF.scala 166:28 167:17 39:22]
  wire [38:0] _GEN_28 = 2'h3 == state ? specialNPCR : 39'h0; // @[NaiveIBF.scala 162:17 98:18]
  wire  _GEN_29 = 2'h3 == state & io_in_valid; // @[NaiveIBF.scala 164:15 98:18]
  wire [1:0] _GEN_31 = 2'h3 == state ? _GEN_26 : state; // @[NaiveIBF.scala 98:18 39:22]
  wire [38:0] _GEN_33 = 2'h2 == state ? _T_148 : _GEN_28; // @[NaiveIBF.scala 150:17 98:18]
  wire  _GEN_34 = 2'h2 == state ? io_in_valid : _GEN_29; // @[NaiveIBF.scala 152:15 98:18]
  wire  _GEN_35 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[NaiveIBF.scala 153:15 98:18]
  wire [1:0] _GEN_36 = 2'h2 == state ? _GEN_24 : _GEN_31; // @[NaiveIBF.scala 98:18]
  wire [2:0] _GEN_37 = 2'h2 == state ? _GEN_25 : pcOffsetR; // @[NaiveIBF.scala 98:18 40:26]
  wire  _GEN_38 = 2'h1 == state ? _T_104 : _GEN_34; // @[NaiveIBF.scala 124:15 98:18]
  wire  _GEN_39 = 2'h1 == state ? _T_105 : _GEN_35; // @[NaiveIBF.scala 125:15 98:18]
  wire [38:0] _GEN_41 = 2'h1 == state ? _T_134 : _GEN_33; // @[NaiveIBF.scala 127:17 98:18]
  wire  canGo = 2'h0 == state ? rvcFinish | rvcNext : _GEN_38; // @[NaiveIBF.scala 100:15 98:18]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[NaiveIBF.scala 101:15 98:18]
  wire [38:0] pnpcOut = 2'h0 == state ? _T_111 : _GEN_41; // @[NaiveIBF.scala 103:17 98:18]
  wire  _T_162 = pnpcOut == _T_132 & _T_4 | pnpcOut == _T_130 & isRVC ? 1'h0 : 1'h1; // @[NaiveIBF.scala 185:27]
  wire  _T_171 = _T_82 | _T_81; // @[NaiveIBF.scala 191:133]
  assign io_in_ready = ~io_in_valid | _T_112 & canIn | loadNextInstline; // @[NaiveIBF.scala 188:60]
  assign io_out_valid = io_in_valid & canGo; // @[NaiveIBF.scala 187:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[NaiveIBF.scala 184:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[NaiveIBF.scala 102:15 98:18]
  assign io_out_bits_pnpc = 2'h0 == state ? _T_111 : _GEN_41; // @[NaiveIBF.scala 103:17 98:18]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_T_82 | _T_81); // @[NaiveIBF.scala 191:87]
  assign io_out_bits_brIdx = {{3'd0}, _T_162}; // @[NaiveIBF.scala 185:21]
  assign io_out_bits_crossPageIPFFix = io_in_bits_exceptionVec_12 & _T_171 & ~specialIPFR; // @[NaiveIBF.scala 192:130]
  always @(posedge clock) begin
    if (reset) begin // @[NaiveIBF.scala 39:22]
      state <= 2'h0; // @[NaiveIBF.scala 39:22]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else begin
        state <= _GEN_36;
      end
    end else begin
      state <= 2'h0; // @[NaiveIBF.scala 172:11]
    end
    if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 40:26]
      pcOffsetR <= 3'h0; // @[NaiveIBF.scala 40:26]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end
    end
    if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 67:28]
      specialIPFR <= 1'h0; // @[NaiveIBF.scala 67:28]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialIPFR <= _GEN_11;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialIPFR <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~flushIFU | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~flushIFU | reset)) begin
          $fatal; // @[NaiveIBF.scala 59:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  specialIPFR = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder(
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_in_bits_crossPageIPFFix,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output [4:0]  io_out_bits_cf_instrType,
  output        io_out_bits_ctrl_src1Type,
  output        io_out_bits_ctrl_src2Type,
  output [3:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output [2:0]  io_out_bits_ctrl_funct3,
  output        io_out_bits_ctrl_func24,
  output        io_out_bits_ctrl_func23,
  output [4:0]  io_out_bits_ctrl_rfSrc1,
  output [4:0]  io_out_bits_ctrl_rfSrc2,
  output [4:0]  io_out_bits_ctrl_rfSrc3,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output        io_out_bits_ctrl_isMou,
  output [63:0] io_out_bits_data_imm,
  output        io_isBranch,
  input         DTLBENABLE,
  input  [63:0] intrVecIDU
);
  wire [63:0] _T = io_in_bits_instr & 64'h707f; // @[Lookup.scala 31:38]
  wire  _T_1 = 64'h13 == _T; // @[Lookup.scala 31:38]
  wire [63:0] _T_2 = io_in_bits_instr & 64'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 64'h1013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 64'h2013 == _T; // @[Lookup.scala 31:38]
  wire  _T_7 = 64'h3013 == _T; // @[Lookup.scala 31:38]
  wire  _T_9 = 64'h4013 == _T; // @[Lookup.scala 31:38]
  wire  _T_11 = 64'h5013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 64'h6013 == _T; // @[Lookup.scala 31:38]
  wire  _T_15 = 64'h7013 == _T; // @[Lookup.scala 31:38]
  wire  _T_17 = 64'h40005013 == _T_2; // @[Lookup.scala 31:38]
  wire [63:0] _T_18 = io_in_bits_instr & 64'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_19 = 64'h33 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_21 = 64'h1033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_23 = 64'h2033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_25 = 64'h3033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_27 = 64'h4033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_29 = 64'h5033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_31 = 64'h6033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_33 = 64'h7033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_35 = 64'h40000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_37 = 64'h40005033 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_38 = io_in_bits_instr & 64'h7f; // @[Lookup.scala 31:38]
  wire  _T_39 = 64'h17 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_41 = 64'h37 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_43 = 64'h6f == _T_38; // @[Lookup.scala 31:38]
  wire  _T_45 = 64'h67 == _T; // @[Lookup.scala 31:38]
  wire  _T_47 = 64'h63 == _T; // @[Lookup.scala 31:38]
  wire  _T_49 = 64'h1063 == _T; // @[Lookup.scala 31:38]
  wire  _T_51 = 64'h4063 == _T; // @[Lookup.scala 31:38]
  wire  _T_53 = 64'h5063 == _T; // @[Lookup.scala 31:38]
  wire  _T_55 = 64'h6063 == _T; // @[Lookup.scala 31:38]
  wire  _T_57 = 64'h7063 == _T; // @[Lookup.scala 31:38]
  wire  _T_59 = 64'h3 == _T; // @[Lookup.scala 31:38]
  wire  _T_61 = 64'h1003 == _T; // @[Lookup.scala 31:38]
  wire  _T_63 = 64'h2003 == _T; // @[Lookup.scala 31:38]
  wire  _T_65 = 64'h4003 == _T; // @[Lookup.scala 31:38]
  wire  _T_67 = 64'h5003 == _T; // @[Lookup.scala 31:38]
  wire  _T_69 = 64'h23 == _T; // @[Lookup.scala 31:38]
  wire  _T_71 = 64'h1023 == _T; // @[Lookup.scala 31:38]
  wire  _T_73 = 64'h2023 == _T; // @[Lookup.scala 31:38]
  wire  _T_75 = 64'h1b == _T; // @[Lookup.scala 31:38]
  wire  _T_77 = 64'h101b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_79 = 64'h501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_81 = 64'h4000501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_83 = 64'h103b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_85 = 64'h503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_87 = 64'h4000503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_89 = 64'h3b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_91 = 64'h4000003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_93 = 64'h6003 == _T; // @[Lookup.scala 31:38]
  wire  _T_95 = 64'h3003 == _T; // @[Lookup.scala 31:38]
  wire  _T_97 = 64'h3023 == _T; // @[Lookup.scala 31:38]
  wire  _T_99 = 64'h6b == _T; // @[Lookup.scala 31:38]
  wire  _T_101 = 64'h2000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_103 = 64'h2001033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_105 = 64'h2002033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_107 = 64'h2003033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_109 = 64'h2004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_111 = 64'h2005033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_113 = 64'h2006033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_115 = 64'h2007033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_117 = 64'h200003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_119 = 64'h200403b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_121 = 64'h200503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_123 = 64'h200603b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_125 = 64'h200703b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_126 = io_in_bits_instr & 64'hffffffff; // @[Lookup.scala 31:38]
  wire  _T_127 = 64'h0 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_128 = io_in_bits_instr & 64'he003; // @[Lookup.scala 31:38]
  wire  _T_129 = 64'h0 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 64'h4000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_133 = 64'h6000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_135 = 64'hc000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_137 = 64'he000 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_138 = io_in_bits_instr & 64'hef83; // @[Lookup.scala 31:38]
  wire  _T_139 = 64'h1 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_141 = 64'h1 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_143 = 64'h2001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_145 = 64'h4001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_147 = 64'h6101 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_149 = 64'h6001 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_150 = io_in_bits_instr & 64'hec03; // @[Lookup.scala 31:38]
  wire  _T_151 = 64'h8001 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_153 = 64'h8401 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_155 = 64'h8801 == _T_150; // @[Lookup.scala 31:38]
  wire [63:0] _T_156 = io_in_bits_instr & 64'hfc63; // @[Lookup.scala 31:38]
  wire  _T_157 = 64'h8c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_159 = 64'h8c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_161 = 64'h8c41 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_163 = 64'h8c61 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_165 = 64'h9c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_167 = 64'h9c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_169 = 64'ha001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_171 = 64'hc001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_173 = 64'he001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_175 = 64'h2 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_177 = 64'h4002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_179 = 64'h6002 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_180 = io_in_bits_instr & 64'hf07f; // @[Lookup.scala 31:38]
  wire  _T_181 = 64'h8002 == _T_180; // @[Lookup.scala 31:38]
  wire [63:0] _T_182 = io_in_bits_instr & 64'hf003; // @[Lookup.scala 31:38]
  wire  _T_183 = 64'h8002 == _T_182; // @[Lookup.scala 31:38]
  wire [63:0] _T_184 = io_in_bits_instr & 64'hffff; // @[Lookup.scala 31:38]
  wire  _T_185 = 64'h9002 == _T_184; // @[Lookup.scala 31:38]
  wire  _T_187 = 64'h9002 == _T_180; // @[Lookup.scala 31:38]
  wire  _T_189 = 64'h9002 == _T_182; // @[Lookup.scala 31:38]
  wire  _T_191 = 64'hc002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_193 = 64'he002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_195 = 64'h73 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_197 = 64'h100073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_199 = 64'h30200073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_201 = 64'hf == _T; // @[Lookup.scala 31:38]
  wire  _T_203 = 64'h10500073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_205 = 64'h10200073 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_206 = io_in_bits_instr & 64'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_207 = 64'h12000073 == _T_206; // @[Lookup.scala 31:38]
  wire [63:0] _T_208 = io_in_bits_instr & 64'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _T_209 = 64'h1000302f == _T_208; // @[Lookup.scala 31:38]
  wire  _T_211 = 64'h1000202f == _T_208; // @[Lookup.scala 31:38]
  wire [63:0] _T_212 = io_in_bits_instr & 64'hf800707f; // @[Lookup.scala 31:38]
  wire  _T_213 = 64'h1800302f == _T_212; // @[Lookup.scala 31:38]
  wire  _T_215 = 64'h1800202f == _T_212; // @[Lookup.scala 31:38]
  wire [63:0] _T_216 = io_in_bits_instr & 64'hf800607f; // @[Lookup.scala 31:38]
  wire  _T_217 = 64'h800202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_219 = 64'h202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_221 = 64'h2000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_223 = 64'h6000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_225 = 64'h4000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_227 = 64'h8000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_229 = 64'ha000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_231 = 64'hc000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_233 = 64'he000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_235 = 64'h1073 == _T; // @[Lookup.scala 31:38]
  wire  _T_237 = 64'h2073 == _T; // @[Lookup.scala 31:38]
  wire  _T_239 = 64'h3073 == _T; // @[Lookup.scala 31:38]
  wire  _T_241 = 64'h5073 == _T; // @[Lookup.scala 31:38]
  wire  _T_243 = 64'h6073 == _T; // @[Lookup.scala 31:38]
  wire  _T_245 = 64'h7073 == _T; // @[Lookup.scala 31:38]
  wire  _T_247 = 64'h100f == _T_126; // @[Lookup.scala 31:38]
  wire  _T_249 = 64'h40000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_251 = 64'h77 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_253 = 64'h10000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_255 = 64'h20000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_257 = 64'h30000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_259 = 64'h42000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_261 = 64'h2000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_263 = 64'h12000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_265 = 64'h22000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_267 = 64'h32000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_269 = 64'h48000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_271 = 64'h8000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_273 = 64'h18000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_275 = 64'h28000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_277 = 64'h38000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_279 = 64'h4a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_281 = 64'ha000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_283 = 64'h1a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_285 = 64'h2a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_287 = 64'h3a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_289 = 64'h44000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_291 = 64'h4000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_293 = 64'h14000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_295 = 64'h24000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_297 = 64'h34000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_299 = 64'h46000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_301 = 64'h6000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_303 = 64'h16000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_305 = 64'h26000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_307 = 64'h36000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_309 = 64'h40002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_311 = 64'h2077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_313 = 64'h10002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_315 = 64'h20002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_317 = 64'h30002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_319 = 64'h42002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_321 = 64'h2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_323 = 64'h12002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_325 = 64'h22002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_327 = 64'h32002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_329 = 64'h44002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_331 = 64'h4002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_333 = 64'h14002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_335 = 64'h24002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_337 = 64'h34002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_339 = 64'h46002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_341 = 64'h6002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_343 = 64'h16002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_345 = 64'h26002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_347 = 64'h36002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_349 = 64'h50000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_351 = 64'h60000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_353 = 64'h52000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_355 = 64'h62000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_357 = 64'h54000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_359 = 64'h64000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_361 = 64'h56000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_363 = 64'h66000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_365 = 64'h58000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_367 = 64'h68000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_369 = 64'h5a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_371 = 64'h6a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_373 = 64'h5c000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_375 = 64'h6c000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_377 = 64'h5e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_379 = 64'h6e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_381 = 64'h50002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_383 = 64'h60002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_385 = 64'h52002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_387 = 64'h62002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_389 = 64'h54002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_391 = 64'h64002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_393 = 64'h56002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_395 = 64'h66002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_397 = 64'h4c000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_399 = 64'hc000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_401 = 64'h1c000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_403 = 64'h2c000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_405 = 64'h3c000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_407 = 64'h4e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_409 = 64'he000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_411 = 64'h1e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_413 = 64'h2e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_415 = 64'h3e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_417 = 64'h80000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_419 = 64'h82000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_421 = 64'h90000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_423 = 64'h92000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_425 = 64'h88000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_427 = 64'h8a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_429 = 64'h98000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_431 = 64'h9a000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_433 = 64'he001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_435 = 64'h1e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_437 = 64'h2e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_439 = 64'h3e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_441 = 64'hfc000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_443 = 64'hfe000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_445 = 64'h80001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_447 = 64'h90001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_449 = 64'ha0001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_451 = 64'hb0001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_453 = 64'h82001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_455 = 64'h92001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_457 = 64'ha2001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_459 = 64'hb2001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_461 = 64'h4001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_463 = 64'h14001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_465 = 64'h6001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_467 = 64'h16001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_469 = 64'h1077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_471 = 64'h10001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_473 = 64'h2001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_475 = 64'h12001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_477 = 64'h6e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_479 = 64'h7e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_481 = 64'h26001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_483 = 64'h20001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_485 = 64'h30001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_487 = 64'h22001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_489 = 64'h32001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_491 = 64'he0000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_493 = 64'h24001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_495 = 64'he6000077 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_496 = io_in_bits_instr & 64'h600707f; // @[Lookup.scala 31:38]
  wire  _T_497 = 64'h6001033 == _T_496; // @[Lookup.scala 31:38]
  wire  _T_499 = 64'hce000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_501 = 64'hf0002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_503 = 64'hb0002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_505 = 64'hc0002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_507 = 64'hd0002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_509 = 64'he0002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_511 = 64'hf2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_513 = 64'hb2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_515 = 64'hc2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_517 = 64'hd2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_519 = 64'he2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_521 = 64'hf4002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_523 = 64'hb4002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_525 = 64'hc4002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_527 = 64'hd4002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_529 = 64'he4002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_531 = 64'hf6002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_533 = 64'hb6002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_535 = 64'hc6002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_537 = 64'hd6002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_539 = 64'he6002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_541 = 64'h90002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_543 = 64'h92002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_545 = 64'ha0002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_547 = 64'ha2002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_549 = 64'h1e002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_551 = 64'h3e002077 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_552 = io_in_bits_instr & 64'hff00707f; // @[Lookup.scala 31:38]
  wire  _T_553 = 64'h70000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_555 = 64'h71000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_557 = 64'h72000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_559 = 64'h73000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_561 = 64'h74000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_563 = 64'h75000077 == _T_552; // @[Lookup.scala 31:38]
  wire [63:0] _T_564 = io_in_bits_instr & 64'hff80707f; // @[Lookup.scala 31:38]
  wire  _T_565 = 64'h78000077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_567 = 64'h78800077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_569 = 64'h7a000077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_571 = 64'h7a800077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_573 = 64'h7c000077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_575 = 64'h7c800077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_577 = 64'h70002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_579 = 64'h80002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_581 = 64'h72002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_583 = 64'h82002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_585 = 64'h74002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_587 = 64'h84002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_589 = 64'h84000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_591 = 64'h85000077 == _T_552; // @[Lookup.scala 31:38]
  wire  _T_593 = 64'h8c000077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_595 = 64'h8d000077 == _T_564; // @[Lookup.scala 31:38]
  wire [63:0] _T_596 = io_in_bits_instr & 64'hfff0707f; // @[Lookup.scala 31:38]
  wire  _T_597 = 64'had100077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_599 = 64'had000077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_601 = 64'had200077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_603 = 64'had400077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_605 = 64'hae800077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_607 = 64'hae900077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_609 = 64'hae000077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_611 = 64'hae100077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_613 = 64'had800077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_615 = 64'hac800077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_617 = 64'hac900077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_619 = 64'haca00077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_621 = 64'hacb00077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_623 = 64'had300077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_625 = 64'hacc00077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_627 = 64'hacd00077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_629 = 64'hace00077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_631 = 64'hacf00077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_633 = 64'had700077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_635 = 64'he4000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_637 = 64'hf4000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_639 = 64'haf800077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_641 = 64'haf900077 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_643 = 64'h36001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_645 = 64'hd4001077 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_647 = 64'he8000077 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_649 = 64'hde000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_651 = 64'hac000077 == _T_564; // @[Lookup.scala 31:38]
  wire  _T_653 = 64'h34001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_655 = 64'ha0000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_657 = 64'hb0000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_659 = 64'ha2000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_661 = 64'hb2000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_663 = 64'h86000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_665 = 64'h96000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_667 = 64'ha8000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_669 = 64'hb8000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_671 = 64'haa000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_673 = 64'hba000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_675 = 64'h8e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_677 = 64'h9e000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_679 = 64'h40001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_681 = 64'h50001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_683 = 64'h62001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_685 = 64'h72001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_687 = 64'h44001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_689 = 64'h54001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_691 = 64'h64001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_693 = 64'h74001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_695 = 64'h8e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_697 = 64'h9e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_699 = 64'hae001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_701 = 64'hbe001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_703 = 64'h8001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_705 = 64'h18001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_707 = 64'h28001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_709 = 64'h38001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_711 = 64'h3a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_713 = 64'h58001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_715 = 64'h68001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_717 = 64'h78001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_719 = 64'h5e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_721 = 64'hc001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_723 = 64'h1c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_725 = 64'h2c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_727 = 64'ha001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_729 = 64'h1a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_731 = 64'h2a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_733 = 64'hf0001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_735 = 64'he0001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_737 = 64'hdc001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_739 = 64'hec001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_741 = 64'hfc001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_743 = 64'hda001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_745 = 64'hea001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_747 = 64'hfa001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_749 = 64'h18002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_751 = 64'h28002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_753 = 64'h38002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_755 = 64'h3a002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_757 = 64'h58002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_759 = 64'h68002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_761 = 64'h78002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_763 = 64'h68805013 == _T_596; // @[Lookup.scala 31:38]
  wire  _T_765 = 64'ha006033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_767 = 64'ha004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_769 = 64'h8004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_771 = 64'h48004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_773 = 64'h400503b == _T_496; // @[Lookup.scala 31:38]
  wire [63:0] _T_774 = io_in_bits_instr & 64'hfdf0707f; // @[Lookup.scala 31:38]
  wire  _T_775 = 64'h69f05013 == _T_774; // @[Lookup.scala 31:38]
  wire  _T_777 = 64'h60001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_779 = 64'h70001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_781 = 64'h42001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_783 = 64'h52001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_785 = 64'h46001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_787 = 64'h56001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_789 = 64'h66001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_791 = 64'h76001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_793 = 64'hce001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_795 = 64'hde001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_797 = 64'hee001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_799 = 64'hfe001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_801 = 64'h5a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_803 = 64'h6a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_805 = 64'h7a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_807 = 64'h48001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_809 = 64'h4a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_811 = 64'h5c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_813 = 64'h6c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_815 = 64'h7c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_817 = 64'h4c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_819 = 64'h4e001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_821 = 64'hc8000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_823 = 64'hca000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_825 = 64'hcc000077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_827 = 64'h84001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_829 = 64'h94001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_831 = 64'ha4001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_833 = 64'hb4001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_835 = 64'h86001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_837 = 64'h96001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_839 = 64'ha6001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_841 = 64'hb6001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_843 = 64'h88001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_845 = 64'h98001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_847 = 64'ha8001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_849 = 64'h8a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_851 = 64'h9a001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_853 = 64'haa001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_855 = 64'h8c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_857 = 64'h9c001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_859 = 64'hac001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_861 = 64'hbc001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_863 = 64'hd2001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_865 = 64'he2001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_867 = 64'hf2001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_869 = 64'hc4001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_871 = 64'hc6001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_873 = 64'hd8001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_875 = 64'he8001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_877 = 64'hf8001077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_879 = 64'h5a002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_881 = 64'h6a002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_883 = 64'h7a002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_885 = 64'h4a002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_887 = 64'h4c002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_889 = 64'h4e002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_891 = 64'h5c002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_893 = 64'h6c002077 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_895 = 64'h7c002077 == _T_18; // @[Lookup.scala 31:38]
  wire [4:0] _T_896 = _T_895 ? 5'h1c : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_897 = _T_893 ? 5'h1c : _T_896; // @[Lookup.scala 33:37]
  wire [4:0] _T_898 = _T_891 ? 5'h1c : _T_897; // @[Lookup.scala 33:37]
  wire [4:0] _T_899 = _T_889 ? 5'h1c : _T_898; // @[Lookup.scala 33:37]
  wire [4:0] _T_900 = _T_887 ? 5'h1c : _T_899; // @[Lookup.scala 33:37]
  wire [4:0] _T_901 = _T_885 ? 5'h1c : _T_900; // @[Lookup.scala 33:37]
  wire [4:0] _T_902 = _T_883 ? 5'h1c : _T_901; // @[Lookup.scala 33:37]
  wire [4:0] _T_903 = _T_881 ? 5'h1c : _T_902; // @[Lookup.scala 33:37]
  wire [4:0] _T_904 = _T_879 ? 5'h1c : _T_903; // @[Lookup.scala 33:37]
  wire [4:0] _T_905 = _T_877 ? 5'h1c : _T_904; // @[Lookup.scala 33:37]
  wire [4:0] _T_906 = _T_875 ? 5'h1c : _T_905; // @[Lookup.scala 33:37]
  wire [4:0] _T_907 = _T_873 ? 5'h1c : _T_906; // @[Lookup.scala 33:37]
  wire [4:0] _T_908 = _T_871 ? 5'h1c : _T_907; // @[Lookup.scala 33:37]
  wire [4:0] _T_909 = _T_869 ? 5'h1c : _T_908; // @[Lookup.scala 33:37]
  wire [4:0] _T_910 = _T_867 ? 5'h1c : _T_909; // @[Lookup.scala 33:37]
  wire [4:0] _T_911 = _T_865 ? 5'h1c : _T_910; // @[Lookup.scala 33:37]
  wire [4:0] _T_912 = _T_863 ? 5'h1c : _T_911; // @[Lookup.scala 33:37]
  wire [4:0] _T_913 = _T_861 ? 5'h1c : _T_912; // @[Lookup.scala 33:37]
  wire [4:0] _T_914 = _T_859 ? 5'h1c : _T_913; // @[Lookup.scala 33:37]
  wire [4:0] _T_915 = _T_857 ? 5'h1c : _T_914; // @[Lookup.scala 33:37]
  wire [4:0] _T_916 = _T_855 ? 5'h1c : _T_915; // @[Lookup.scala 33:37]
  wire [4:0] _T_917 = _T_853 ? 5'h1c : _T_916; // @[Lookup.scala 33:37]
  wire [4:0] _T_918 = _T_851 ? 5'h1c : _T_917; // @[Lookup.scala 33:37]
  wire [4:0] _T_919 = _T_849 ? 5'h1c : _T_918; // @[Lookup.scala 33:37]
  wire [4:0] _T_920 = _T_847 ? 5'h1c : _T_919; // @[Lookup.scala 33:37]
  wire [4:0] _T_921 = _T_845 ? 5'h1c : _T_920; // @[Lookup.scala 33:37]
  wire [4:0] _T_922 = _T_843 ? 5'h1c : _T_921; // @[Lookup.scala 33:37]
  wire [4:0] _T_923 = _T_841 ? 5'h1c : _T_922; // @[Lookup.scala 33:37]
  wire [4:0] _T_924 = _T_839 ? 5'h1c : _T_923; // @[Lookup.scala 33:37]
  wire [4:0] _T_925 = _T_837 ? 5'h1c : _T_924; // @[Lookup.scala 33:37]
  wire [4:0] _T_926 = _T_835 ? 5'h1c : _T_925; // @[Lookup.scala 33:37]
  wire [4:0] _T_927 = _T_833 ? 5'h1c : _T_926; // @[Lookup.scala 33:37]
  wire [4:0] _T_928 = _T_831 ? 5'h1c : _T_927; // @[Lookup.scala 33:37]
  wire [4:0] _T_929 = _T_829 ? 5'h1c : _T_928; // @[Lookup.scala 33:37]
  wire [4:0] _T_930 = _T_827 ? 5'h1c : _T_929; // @[Lookup.scala 33:37]
  wire [4:0] _T_931 = _T_825 ? 5'h1c : _T_930; // @[Lookup.scala 33:37]
  wire [4:0] _T_932 = _T_823 ? 5'h1c : _T_931; // @[Lookup.scala 33:37]
  wire [4:0] _T_933 = _T_821 ? 5'h1c : _T_932; // @[Lookup.scala 33:37]
  wire [4:0] _T_934 = _T_819 ? 5'h1c : _T_933; // @[Lookup.scala 33:37]
  wire [4:0] _T_935 = _T_817 ? 5'h1c : _T_934; // @[Lookup.scala 33:37]
  wire [4:0] _T_936 = _T_815 ? 5'h1c : _T_935; // @[Lookup.scala 33:37]
  wire [4:0] _T_937 = _T_813 ? 5'h1c : _T_936; // @[Lookup.scala 33:37]
  wire [4:0] _T_938 = _T_811 ? 5'h1c : _T_937; // @[Lookup.scala 33:37]
  wire [4:0] _T_939 = _T_809 ? 5'h1c : _T_938; // @[Lookup.scala 33:37]
  wire [4:0] _T_940 = _T_807 ? 5'h1c : _T_939; // @[Lookup.scala 33:37]
  wire [4:0] _T_941 = _T_805 ? 5'h1c : _T_940; // @[Lookup.scala 33:37]
  wire [4:0] _T_942 = _T_803 ? 5'h1c : _T_941; // @[Lookup.scala 33:37]
  wire [4:0] _T_943 = _T_801 ? 5'h1c : _T_942; // @[Lookup.scala 33:37]
  wire [4:0] _T_944 = _T_799 ? 5'h1c : _T_943; // @[Lookup.scala 33:37]
  wire [4:0] _T_945 = _T_797 ? 5'h1c : _T_944; // @[Lookup.scala 33:37]
  wire [4:0] _T_946 = _T_795 ? 5'h1c : _T_945; // @[Lookup.scala 33:37]
  wire [4:0] _T_947 = _T_793 ? 5'h1c : _T_946; // @[Lookup.scala 33:37]
  wire [4:0] _T_948 = _T_791 ? 5'h1c : _T_947; // @[Lookup.scala 33:37]
  wire [4:0] _T_949 = _T_789 ? 5'h1c : _T_948; // @[Lookup.scala 33:37]
  wire [4:0] _T_950 = _T_787 ? 5'h1c : _T_949; // @[Lookup.scala 33:37]
  wire [4:0] _T_951 = _T_785 ? 5'h1c : _T_950; // @[Lookup.scala 33:37]
  wire [4:0] _T_952 = _T_783 ? 5'h1c : _T_951; // @[Lookup.scala 33:37]
  wire [4:0] _T_953 = _T_781 ? 5'h1c : _T_952; // @[Lookup.scala 33:37]
  wire [4:0] _T_954 = _T_779 ? 5'h1c : _T_953; // @[Lookup.scala 33:37]
  wire [4:0] _T_955 = _T_777 ? 5'h1c : _T_954; // @[Lookup.scala 33:37]
  wire [4:0] _T_956 = _T_775 ? 5'h17 : _T_955; // @[Lookup.scala 33:37]
  wire [4:0] _T_957 = _T_773 ? 5'h14 : _T_956; // @[Lookup.scala 33:37]
  wire [4:0] _T_958 = _T_771 ? 5'h14 : _T_957; // @[Lookup.scala 33:37]
  wire [4:0] _T_959 = _T_769 ? 5'h14 : _T_958; // @[Lookup.scala 33:37]
  wire [4:0] _T_960 = _T_767 ? 5'h14 : _T_959; // @[Lookup.scala 33:37]
  wire [4:0] _T_961 = _T_765 ? 5'h14 : _T_960; // @[Lookup.scala 33:37]
  wire [4:0] _T_962 = _T_763 ? 5'h17 : _T_961; // @[Lookup.scala 33:37]
  wire [4:0] _T_963 = _T_761 ? 5'h16 : _T_962; // @[Lookup.scala 33:37]
  wire [4:0] _T_964 = _T_759 ? 5'h16 : _T_963; // @[Lookup.scala 33:37]
  wire [4:0] _T_965 = _T_757 ? 5'h16 : _T_964; // @[Lookup.scala 33:37]
  wire [4:0] _T_966 = _T_755 ? 5'h16 : _T_965; // @[Lookup.scala 33:37]
  wire [4:0] _T_967 = _T_753 ? 5'h16 : _T_966; // @[Lookup.scala 33:37]
  wire [4:0] _T_968 = _T_751 ? 5'h16 : _T_967; // @[Lookup.scala 33:37]
  wire [4:0] _T_969 = _T_749 ? 5'h16 : _T_968; // @[Lookup.scala 33:37]
  wire [4:0] _T_970 = _T_747 ? 5'h16 : _T_969; // @[Lookup.scala 33:37]
  wire [4:0] _T_971 = _T_745 ? 5'h16 : _T_970; // @[Lookup.scala 33:37]
  wire [4:0] _T_972 = _T_743 ? 5'h16 : _T_971; // @[Lookup.scala 33:37]
  wire [4:0] _T_973 = _T_741 ? 5'h16 : _T_972; // @[Lookup.scala 33:37]
  wire [4:0] _T_974 = _T_739 ? 5'h16 : _T_973; // @[Lookup.scala 33:37]
  wire [4:0] _T_975 = _T_737 ? 5'h16 : _T_974; // @[Lookup.scala 33:37]
  wire [4:0] _T_976 = _T_735 ? 5'h16 : _T_975; // @[Lookup.scala 33:37]
  wire [4:0] _T_977 = _T_733 ? 5'h16 : _T_976; // @[Lookup.scala 33:37]
  wire [4:0] _T_978 = _T_731 ? 5'h16 : _T_977; // @[Lookup.scala 33:37]
  wire [4:0] _T_979 = _T_729 ? 5'h16 : _T_978; // @[Lookup.scala 33:37]
  wire [4:0] _T_980 = _T_727 ? 5'h16 : _T_979; // @[Lookup.scala 33:37]
  wire [4:0] _T_981 = _T_725 ? 5'h16 : _T_980; // @[Lookup.scala 33:37]
  wire [4:0] _T_982 = _T_723 ? 5'h16 : _T_981; // @[Lookup.scala 33:37]
  wire [4:0] _T_983 = _T_721 ? 5'h16 : _T_982; // @[Lookup.scala 33:37]
  wire [4:0] _T_984 = _T_719 ? 5'h16 : _T_983; // @[Lookup.scala 33:37]
  wire [4:0] _T_985 = _T_717 ? 5'h16 : _T_984; // @[Lookup.scala 33:37]
  wire [4:0] _T_986 = _T_715 ? 5'h16 : _T_985; // @[Lookup.scala 33:37]
  wire [4:0] _T_987 = _T_713 ? 5'h16 : _T_986; // @[Lookup.scala 33:37]
  wire [4:0] _T_988 = _T_711 ? 5'h16 : _T_987; // @[Lookup.scala 33:37]
  wire [4:0] _T_989 = _T_709 ? 5'h16 : _T_988; // @[Lookup.scala 33:37]
  wire [4:0] _T_990 = _T_707 ? 5'h16 : _T_989; // @[Lookup.scala 33:37]
  wire [4:0] _T_991 = _T_705 ? 5'h16 : _T_990; // @[Lookup.scala 33:37]
  wire [4:0] _T_992 = _T_703 ? 5'h16 : _T_991; // @[Lookup.scala 33:37]
  wire [4:0] _T_993 = _T_701 ? 5'h16 : _T_992; // @[Lookup.scala 33:37]
  wire [4:0] _T_994 = _T_699 ? 5'h16 : _T_993; // @[Lookup.scala 33:37]
  wire [4:0] _T_995 = _T_697 ? 5'h16 : _T_994; // @[Lookup.scala 33:37]
  wire [4:0] _T_996 = _T_695 ? 5'h16 : _T_995; // @[Lookup.scala 33:37]
  wire [4:0] _T_997 = _T_693 ? 5'h16 : _T_996; // @[Lookup.scala 33:37]
  wire [4:0] _T_998 = _T_691 ? 5'h16 : _T_997; // @[Lookup.scala 33:37]
  wire [4:0] _T_999 = _T_689 ? 5'h16 : _T_998; // @[Lookup.scala 33:37]
  wire [4:0] _T_1000 = _T_687 ? 5'h16 : _T_999; // @[Lookup.scala 33:37]
  wire [4:0] _T_1001 = _T_685 ? 5'h16 : _T_1000; // @[Lookup.scala 33:37]
  wire [4:0] _T_1002 = _T_683 ? 5'h16 : _T_1001; // @[Lookup.scala 33:37]
  wire [4:0] _T_1003 = _T_681 ? 5'h16 : _T_1002; // @[Lookup.scala 33:37]
  wire [4:0] _T_1004 = _T_679 ? 5'h16 : _T_1003; // @[Lookup.scala 33:37]
  wire [4:0] _T_1005 = _T_677 ? 5'h16 : _T_1004; // @[Lookup.scala 33:37]
  wire [4:0] _T_1006 = _T_675 ? 5'h16 : _T_1005; // @[Lookup.scala 33:37]
  wire [4:0] _T_1007 = _T_673 ? 5'h16 : _T_1006; // @[Lookup.scala 33:37]
  wire [4:0] _T_1008 = _T_671 ? 5'h16 : _T_1007; // @[Lookup.scala 33:37]
  wire [4:0] _T_1009 = _T_669 ? 5'h16 : _T_1008; // @[Lookup.scala 33:37]
  wire [4:0] _T_1010 = _T_667 ? 5'h16 : _T_1009; // @[Lookup.scala 33:37]
  wire [4:0] _T_1011 = _T_665 ? 5'h16 : _T_1010; // @[Lookup.scala 33:37]
  wire [4:0] _T_1012 = _T_663 ? 5'h16 : _T_1011; // @[Lookup.scala 33:37]
  wire [4:0] _T_1013 = _T_661 ? 5'h16 : _T_1012; // @[Lookup.scala 33:37]
  wire [4:0] _T_1014 = _T_659 ? 5'h16 : _T_1013; // @[Lookup.scala 33:37]
  wire [4:0] _T_1015 = _T_657 ? 5'h16 : _T_1014; // @[Lookup.scala 33:37]
  wire [4:0] _T_1016 = _T_655 ? 5'h16 : _T_1015; // @[Lookup.scala 33:37]
  wire [4:0] _T_1017 = _T_653 ? 5'h15 : _T_1016; // @[Lookup.scala 33:37]
  wire [4:0] _T_1018 = _T_651 ? 5'h15 : _T_1017; // @[Lookup.scala 33:37]
  wire [4:0] _T_1019 = _T_649 ? 5'h15 : _T_1018; // @[Lookup.scala 33:37]
  wire [4:0] _T_1020 = _T_647 ? 5'h15 : _T_1019; // @[Lookup.scala 33:37]
  wire [4:0] _T_1021 = _T_645 ? 5'h15 : _T_1020; // @[Lookup.scala 33:37]
  wire [4:0] _T_1022 = _T_643 ? 5'h15 : _T_1021; // @[Lookup.scala 33:37]
  wire [4:0] _T_1023 = _T_641 ? 5'h15 : _T_1022; // @[Lookup.scala 33:37]
  wire [4:0] _T_1024 = _T_639 ? 5'h15 : _T_1023; // @[Lookup.scala 33:37]
  wire [4:0] _T_1025 = _T_637 ? 5'h15 : _T_1024; // @[Lookup.scala 33:37]
  wire [4:0] _T_1026 = _T_635 ? 5'h15 : _T_1025; // @[Lookup.scala 33:37]
  wire [4:0] _T_1027 = _T_633 ? 5'h15 : _T_1026; // @[Lookup.scala 33:37]
  wire [4:0] _T_1028 = _T_631 ? 5'h15 : _T_1027; // @[Lookup.scala 33:37]
  wire [4:0] _T_1029 = _T_629 ? 5'h15 : _T_1028; // @[Lookup.scala 33:37]
  wire [4:0] _T_1030 = _T_627 ? 5'h15 : _T_1029; // @[Lookup.scala 33:37]
  wire [4:0] _T_1031 = _T_625 ? 5'h15 : _T_1030; // @[Lookup.scala 33:37]
  wire [4:0] _T_1032 = _T_623 ? 5'h15 : _T_1031; // @[Lookup.scala 33:37]
  wire [4:0] _T_1033 = _T_621 ? 5'h15 : _T_1032; // @[Lookup.scala 33:37]
  wire [4:0] _T_1034 = _T_619 ? 5'h15 : _T_1033; // @[Lookup.scala 33:37]
  wire [4:0] _T_1035 = _T_617 ? 5'h15 : _T_1034; // @[Lookup.scala 33:37]
  wire [4:0] _T_1036 = _T_615 ? 5'h15 : _T_1035; // @[Lookup.scala 33:37]
  wire [4:0] _T_1037 = _T_613 ? 5'h15 : _T_1036; // @[Lookup.scala 33:37]
  wire [4:0] _T_1038 = _T_611 ? 5'h15 : _T_1037; // @[Lookup.scala 33:37]
  wire [4:0] _T_1039 = _T_609 ? 5'h15 : _T_1038; // @[Lookup.scala 33:37]
  wire [4:0] _T_1040 = _T_607 ? 5'h15 : _T_1039; // @[Lookup.scala 33:37]
  wire [4:0] _T_1041 = _T_605 ? 5'h15 : _T_1040; // @[Lookup.scala 33:37]
  wire [4:0] _T_1042 = _T_603 ? 5'h15 : _T_1041; // @[Lookup.scala 33:37]
  wire [4:0] _T_1043 = _T_601 ? 5'h15 : _T_1042; // @[Lookup.scala 33:37]
  wire [4:0] _T_1044 = _T_599 ? 5'h15 : _T_1043; // @[Lookup.scala 33:37]
  wire [4:0] _T_1045 = _T_597 ? 5'h15 : _T_1044; // @[Lookup.scala 33:37]
  wire [4:0] _T_1046 = _T_595 ? 5'h15 : _T_1045; // @[Lookup.scala 33:37]
  wire [4:0] _T_1047 = _T_593 ? 5'h15 : _T_1046; // @[Lookup.scala 33:37]
  wire [4:0] _T_1048 = _T_591 ? 5'h15 : _T_1047; // @[Lookup.scala 33:37]
  wire [4:0] _T_1049 = _T_589 ? 5'h15 : _T_1048; // @[Lookup.scala 33:37]
  wire [4:0] _T_1050 = _T_587 ? 5'h15 : _T_1049; // @[Lookup.scala 33:37]
  wire [4:0] _T_1051 = _T_585 ? 5'h15 : _T_1050; // @[Lookup.scala 33:37]
  wire [4:0] _T_1052 = _T_583 ? 5'h15 : _T_1051; // @[Lookup.scala 33:37]
  wire [4:0] _T_1053 = _T_581 ? 5'h15 : _T_1052; // @[Lookup.scala 33:37]
  wire [4:0] _T_1054 = _T_579 ? 5'h15 : _T_1053; // @[Lookup.scala 33:37]
  wire [4:0] _T_1055 = _T_577 ? 5'h15 : _T_1054; // @[Lookup.scala 33:37]
  wire [4:0] _T_1056 = _T_575 ? 5'h15 : _T_1055; // @[Lookup.scala 33:37]
  wire [4:0] _T_1057 = _T_573 ? 5'h15 : _T_1056; // @[Lookup.scala 33:37]
  wire [4:0] _T_1058 = _T_571 ? 5'h15 : _T_1057; // @[Lookup.scala 33:37]
  wire [4:0] _T_1059 = _T_569 ? 5'h15 : _T_1058; // @[Lookup.scala 33:37]
  wire [4:0] _T_1060 = _T_567 ? 5'h15 : _T_1059; // @[Lookup.scala 33:37]
  wire [4:0] _T_1061 = _T_565 ? 5'h15 : _T_1060; // @[Lookup.scala 33:37]
  wire [4:0] _T_1062 = _T_563 ? 5'h15 : _T_1061; // @[Lookup.scala 33:37]
  wire [4:0] _T_1063 = _T_561 ? 5'h15 : _T_1062; // @[Lookup.scala 33:37]
  wire [4:0] _T_1064 = _T_559 ? 5'h15 : _T_1063; // @[Lookup.scala 33:37]
  wire [4:0] _T_1065 = _T_557 ? 5'h15 : _T_1064; // @[Lookup.scala 33:37]
  wire [4:0] _T_1066 = _T_555 ? 5'h15 : _T_1065; // @[Lookup.scala 33:37]
  wire [4:0] _T_1067 = _T_553 ? 5'h15 : _T_1066; // @[Lookup.scala 33:37]
  wire [4:0] _T_1068 = _T_551 ? 5'h14 : _T_1067; // @[Lookup.scala 33:37]
  wire [4:0] _T_1069 = _T_549 ? 5'h14 : _T_1068; // @[Lookup.scala 33:37]
  wire [4:0] _T_1070 = _T_547 ? 5'h14 : _T_1069; // @[Lookup.scala 33:37]
  wire [4:0] _T_1071 = _T_545 ? 5'h14 : _T_1070; // @[Lookup.scala 33:37]
  wire [4:0] _T_1072 = _T_543 ? 5'h14 : _T_1071; // @[Lookup.scala 33:37]
  wire [4:0] _T_1073 = _T_541 ? 5'h14 : _T_1072; // @[Lookup.scala 33:37]
  wire [4:0] _T_1074 = _T_539 ? 5'h14 : _T_1073; // @[Lookup.scala 33:37]
  wire [4:0] _T_1075 = _T_537 ? 5'h14 : _T_1074; // @[Lookup.scala 33:37]
  wire [4:0] _T_1076 = _T_535 ? 5'h14 : _T_1075; // @[Lookup.scala 33:37]
  wire [4:0] _T_1077 = _T_533 ? 5'h14 : _T_1076; // @[Lookup.scala 33:37]
  wire [4:0] _T_1078 = _T_531 ? 5'h14 : _T_1077; // @[Lookup.scala 33:37]
  wire [4:0] _T_1079 = _T_529 ? 5'h14 : _T_1078; // @[Lookup.scala 33:37]
  wire [4:0] _T_1080 = _T_527 ? 5'h14 : _T_1079; // @[Lookup.scala 33:37]
  wire [4:0] _T_1081 = _T_525 ? 5'h14 : _T_1080; // @[Lookup.scala 33:37]
  wire [4:0] _T_1082 = _T_523 ? 5'h14 : _T_1081; // @[Lookup.scala 33:37]
  wire [4:0] _T_1083 = _T_521 ? 5'h14 : _T_1082; // @[Lookup.scala 33:37]
  wire [4:0] _T_1084 = _T_519 ? 5'h14 : _T_1083; // @[Lookup.scala 33:37]
  wire [4:0] _T_1085 = _T_517 ? 5'h14 : _T_1084; // @[Lookup.scala 33:37]
  wire [4:0] _T_1086 = _T_515 ? 5'h14 : _T_1085; // @[Lookup.scala 33:37]
  wire [4:0] _T_1087 = _T_513 ? 5'h14 : _T_1086; // @[Lookup.scala 33:37]
  wire [4:0] _T_1088 = _T_511 ? 5'h14 : _T_1087; // @[Lookup.scala 33:37]
  wire [4:0] _T_1089 = _T_509 ? 5'h14 : _T_1088; // @[Lookup.scala 33:37]
  wire [4:0] _T_1090 = _T_507 ? 5'h14 : _T_1089; // @[Lookup.scala 33:37]
  wire [4:0] _T_1091 = _T_505 ? 5'h14 : _T_1090; // @[Lookup.scala 33:37]
  wire [4:0] _T_1092 = _T_503 ? 5'h14 : _T_1091; // @[Lookup.scala 33:37]
  wire [4:0] _T_1093 = _T_501 ? 5'h14 : _T_1092; // @[Lookup.scala 33:37]
  wire [4:0] _T_1094 = _T_499 ? 5'h14 : _T_1093; // @[Lookup.scala 33:37]
  wire [4:0] _T_1095 = _T_497 ? 5'h14 : _T_1094; // @[Lookup.scala 33:37]
  wire [4:0] _T_1096 = _T_495 ? 5'h14 : _T_1095; // @[Lookup.scala 33:37]
  wire [4:0] _T_1097 = _T_493 ? 5'h14 : _T_1096; // @[Lookup.scala 33:37]
  wire [4:0] _T_1098 = _T_491 ? 5'h14 : _T_1097; // @[Lookup.scala 33:37]
  wire [4:0] _T_1099 = _T_489 ? 5'h14 : _T_1098; // @[Lookup.scala 33:37]
  wire [4:0] _T_1100 = _T_487 ? 5'h14 : _T_1099; // @[Lookup.scala 33:37]
  wire [4:0] _T_1101 = _T_485 ? 5'h14 : _T_1100; // @[Lookup.scala 33:37]
  wire [4:0] _T_1102 = _T_483 ? 5'h14 : _T_1101; // @[Lookup.scala 33:37]
  wire [4:0] _T_1103 = _T_481 ? 5'h14 : _T_1102; // @[Lookup.scala 33:37]
  wire [4:0] _T_1104 = _T_479 ? 5'h14 : _T_1103; // @[Lookup.scala 33:37]
  wire [4:0] _T_1105 = _T_477 ? 5'h14 : _T_1104; // @[Lookup.scala 33:37]
  wire [4:0] _T_1106 = _T_475 ? 5'h14 : _T_1105; // @[Lookup.scala 33:37]
  wire [4:0] _T_1107 = _T_473 ? 5'h14 : _T_1106; // @[Lookup.scala 33:37]
  wire [4:0] _T_1108 = _T_471 ? 5'h14 : _T_1107; // @[Lookup.scala 33:37]
  wire [4:0] _T_1109 = _T_469 ? 5'h14 : _T_1108; // @[Lookup.scala 33:37]
  wire [4:0] _T_1110 = _T_467 ? 5'h14 : _T_1109; // @[Lookup.scala 33:37]
  wire [4:0] _T_1111 = _T_465 ? 5'h14 : _T_1110; // @[Lookup.scala 33:37]
  wire [4:0] _T_1112 = _T_463 ? 5'h14 : _T_1111; // @[Lookup.scala 33:37]
  wire [4:0] _T_1113 = _T_461 ? 5'h14 : _T_1112; // @[Lookup.scala 33:37]
  wire [4:0] _T_1114 = _T_459 ? 5'h14 : _T_1113; // @[Lookup.scala 33:37]
  wire [4:0] _T_1115 = _T_457 ? 5'h14 : _T_1114; // @[Lookup.scala 33:37]
  wire [4:0] _T_1116 = _T_455 ? 5'h14 : _T_1115; // @[Lookup.scala 33:37]
  wire [4:0] _T_1117 = _T_453 ? 5'h14 : _T_1116; // @[Lookup.scala 33:37]
  wire [4:0] _T_1118 = _T_451 ? 5'h14 : _T_1117; // @[Lookup.scala 33:37]
  wire [4:0] _T_1119 = _T_449 ? 5'h14 : _T_1118; // @[Lookup.scala 33:37]
  wire [4:0] _T_1120 = _T_447 ? 5'h14 : _T_1119; // @[Lookup.scala 33:37]
  wire [4:0] _T_1121 = _T_445 ? 5'h14 : _T_1120; // @[Lookup.scala 33:37]
  wire [4:0] _T_1122 = _T_443 ? 5'h14 : _T_1121; // @[Lookup.scala 33:37]
  wire [4:0] _T_1123 = _T_441 ? 5'h14 : _T_1122; // @[Lookup.scala 33:37]
  wire [4:0] _T_1124 = _T_439 ? 5'h14 : _T_1123; // @[Lookup.scala 33:37]
  wire [4:0] _T_1125 = _T_437 ? 5'h14 : _T_1124; // @[Lookup.scala 33:37]
  wire [4:0] _T_1126 = _T_435 ? 5'h14 : _T_1125; // @[Lookup.scala 33:37]
  wire [4:0] _T_1127 = _T_433 ? 5'h14 : _T_1126; // @[Lookup.scala 33:37]
  wire [4:0] _T_1128 = _T_431 ? 5'h14 : _T_1127; // @[Lookup.scala 33:37]
  wire [4:0] _T_1129 = _T_429 ? 5'h14 : _T_1128; // @[Lookup.scala 33:37]
  wire [4:0] _T_1130 = _T_427 ? 5'h14 : _T_1129; // @[Lookup.scala 33:37]
  wire [4:0] _T_1131 = _T_425 ? 5'h14 : _T_1130; // @[Lookup.scala 33:37]
  wire [4:0] _T_1132 = _T_423 ? 5'h14 : _T_1131; // @[Lookup.scala 33:37]
  wire [4:0] _T_1133 = _T_421 ? 5'h14 : _T_1132; // @[Lookup.scala 33:37]
  wire [4:0] _T_1134 = _T_419 ? 5'h14 : _T_1133; // @[Lookup.scala 33:37]
  wire [4:0] _T_1135 = _T_417 ? 5'h14 : _T_1134; // @[Lookup.scala 33:37]
  wire [4:0] _T_1136 = _T_415 ? 5'h14 : _T_1135; // @[Lookup.scala 33:37]
  wire [4:0] _T_1137 = _T_413 ? 5'h14 : _T_1136; // @[Lookup.scala 33:37]
  wire [4:0] _T_1138 = _T_411 ? 5'h14 : _T_1137; // @[Lookup.scala 33:37]
  wire [4:0] _T_1139 = _T_409 ? 5'h14 : _T_1138; // @[Lookup.scala 33:37]
  wire [4:0] _T_1140 = _T_407 ? 5'h14 : _T_1139; // @[Lookup.scala 33:37]
  wire [4:0] _T_1141 = _T_405 ? 5'h14 : _T_1140; // @[Lookup.scala 33:37]
  wire [4:0] _T_1142 = _T_403 ? 5'h14 : _T_1141; // @[Lookup.scala 33:37]
  wire [4:0] _T_1143 = _T_401 ? 5'h14 : _T_1142; // @[Lookup.scala 33:37]
  wire [4:0] _T_1144 = _T_399 ? 5'h14 : _T_1143; // @[Lookup.scala 33:37]
  wire [4:0] _T_1145 = _T_397 ? 5'h14 : _T_1144; // @[Lookup.scala 33:37]
  wire [4:0] _T_1146 = _T_395 ? 5'h14 : _T_1145; // @[Lookup.scala 33:37]
  wire [4:0] _T_1147 = _T_393 ? 5'h14 : _T_1146; // @[Lookup.scala 33:37]
  wire [4:0] _T_1148 = _T_391 ? 5'h14 : _T_1147; // @[Lookup.scala 33:37]
  wire [4:0] _T_1149 = _T_389 ? 5'h14 : _T_1148; // @[Lookup.scala 33:37]
  wire [4:0] _T_1150 = _T_387 ? 5'h14 : _T_1149; // @[Lookup.scala 33:37]
  wire [4:0] _T_1151 = _T_385 ? 5'h14 : _T_1150; // @[Lookup.scala 33:37]
  wire [4:0] _T_1152 = _T_383 ? 5'h14 : _T_1151; // @[Lookup.scala 33:37]
  wire [4:0] _T_1153 = _T_381 ? 5'h14 : _T_1152; // @[Lookup.scala 33:37]
  wire [4:0] _T_1154 = _T_379 ? 5'h14 : _T_1153; // @[Lookup.scala 33:37]
  wire [4:0] _T_1155 = _T_377 ? 5'h14 : _T_1154; // @[Lookup.scala 33:37]
  wire [4:0] _T_1156 = _T_375 ? 5'h14 : _T_1155; // @[Lookup.scala 33:37]
  wire [4:0] _T_1157 = _T_373 ? 5'h14 : _T_1156; // @[Lookup.scala 33:37]
  wire [4:0] _T_1158 = _T_371 ? 5'h14 : _T_1157; // @[Lookup.scala 33:37]
  wire [4:0] _T_1159 = _T_369 ? 5'h14 : _T_1158; // @[Lookup.scala 33:37]
  wire [4:0] _T_1160 = _T_367 ? 5'h14 : _T_1159; // @[Lookup.scala 33:37]
  wire [4:0] _T_1161 = _T_365 ? 5'h14 : _T_1160; // @[Lookup.scala 33:37]
  wire [4:0] _T_1162 = _T_363 ? 5'h14 : _T_1161; // @[Lookup.scala 33:37]
  wire [4:0] _T_1163 = _T_361 ? 5'h14 : _T_1162; // @[Lookup.scala 33:37]
  wire [4:0] _T_1164 = _T_359 ? 5'h14 : _T_1163; // @[Lookup.scala 33:37]
  wire [4:0] _T_1165 = _T_357 ? 5'h14 : _T_1164; // @[Lookup.scala 33:37]
  wire [4:0] _T_1166 = _T_355 ? 5'h14 : _T_1165; // @[Lookup.scala 33:37]
  wire [4:0] _T_1167 = _T_353 ? 5'h14 : _T_1166; // @[Lookup.scala 33:37]
  wire [4:0] _T_1168 = _T_351 ? 5'h14 : _T_1167; // @[Lookup.scala 33:37]
  wire [4:0] _T_1169 = _T_349 ? 5'h14 : _T_1168; // @[Lookup.scala 33:37]
  wire [4:0] _T_1170 = _T_347 ? 5'h14 : _T_1169; // @[Lookup.scala 33:37]
  wire [4:0] _T_1171 = _T_345 ? 5'h14 : _T_1170; // @[Lookup.scala 33:37]
  wire [4:0] _T_1172 = _T_343 ? 5'h14 : _T_1171; // @[Lookup.scala 33:37]
  wire [4:0] _T_1173 = _T_341 ? 5'h14 : _T_1172; // @[Lookup.scala 33:37]
  wire [4:0] _T_1174 = _T_339 ? 5'h14 : _T_1173; // @[Lookup.scala 33:37]
  wire [4:0] _T_1175 = _T_337 ? 5'h14 : _T_1174; // @[Lookup.scala 33:37]
  wire [4:0] _T_1176 = _T_335 ? 5'h14 : _T_1175; // @[Lookup.scala 33:37]
  wire [4:0] _T_1177 = _T_333 ? 5'h14 : _T_1176; // @[Lookup.scala 33:37]
  wire [4:0] _T_1178 = _T_331 ? 5'h14 : _T_1177; // @[Lookup.scala 33:37]
  wire [4:0] _T_1179 = _T_329 ? 5'h14 : _T_1178; // @[Lookup.scala 33:37]
  wire [4:0] _T_1180 = _T_327 ? 5'h14 : _T_1179; // @[Lookup.scala 33:37]
  wire [4:0] _T_1181 = _T_325 ? 5'h14 : _T_1180; // @[Lookup.scala 33:37]
  wire [4:0] _T_1182 = _T_323 ? 5'h14 : _T_1181; // @[Lookup.scala 33:37]
  wire [4:0] _T_1183 = _T_321 ? 5'h14 : _T_1182; // @[Lookup.scala 33:37]
  wire [4:0] _T_1184 = _T_319 ? 5'h14 : _T_1183; // @[Lookup.scala 33:37]
  wire [4:0] _T_1185 = _T_317 ? 5'h14 : _T_1184; // @[Lookup.scala 33:37]
  wire [4:0] _T_1186 = _T_315 ? 5'h14 : _T_1185; // @[Lookup.scala 33:37]
  wire [4:0] _T_1187 = _T_313 ? 5'h14 : _T_1186; // @[Lookup.scala 33:37]
  wire [4:0] _T_1188 = _T_311 ? 5'h14 : _T_1187; // @[Lookup.scala 33:37]
  wire [4:0] _T_1189 = _T_309 ? 5'h14 : _T_1188; // @[Lookup.scala 33:37]
  wire [4:0] _T_1190 = _T_307 ? 5'h14 : _T_1189; // @[Lookup.scala 33:37]
  wire [4:0] _T_1191 = _T_305 ? 5'h14 : _T_1190; // @[Lookup.scala 33:37]
  wire [4:0] _T_1192 = _T_303 ? 5'h14 : _T_1191; // @[Lookup.scala 33:37]
  wire [4:0] _T_1193 = _T_301 ? 5'h14 : _T_1192; // @[Lookup.scala 33:37]
  wire [4:0] _T_1194 = _T_299 ? 5'h14 : _T_1193; // @[Lookup.scala 33:37]
  wire [4:0] _T_1195 = _T_297 ? 5'h14 : _T_1194; // @[Lookup.scala 33:37]
  wire [4:0] _T_1196 = _T_295 ? 5'h14 : _T_1195; // @[Lookup.scala 33:37]
  wire [4:0] _T_1197 = _T_293 ? 5'h14 : _T_1196; // @[Lookup.scala 33:37]
  wire [4:0] _T_1198 = _T_291 ? 5'h14 : _T_1197; // @[Lookup.scala 33:37]
  wire [4:0] _T_1199 = _T_289 ? 5'h14 : _T_1198; // @[Lookup.scala 33:37]
  wire [4:0] _T_1200 = _T_287 ? 5'h14 : _T_1199; // @[Lookup.scala 33:37]
  wire [4:0] _T_1201 = _T_285 ? 5'h14 : _T_1200; // @[Lookup.scala 33:37]
  wire [4:0] _T_1202 = _T_283 ? 5'h14 : _T_1201; // @[Lookup.scala 33:37]
  wire [4:0] _T_1203 = _T_281 ? 5'h14 : _T_1202; // @[Lookup.scala 33:37]
  wire [4:0] _T_1204 = _T_279 ? 5'h14 : _T_1203; // @[Lookup.scala 33:37]
  wire [4:0] _T_1205 = _T_277 ? 5'h14 : _T_1204; // @[Lookup.scala 33:37]
  wire [4:0] _T_1206 = _T_275 ? 5'h14 : _T_1205; // @[Lookup.scala 33:37]
  wire [4:0] _T_1207 = _T_273 ? 5'h14 : _T_1206; // @[Lookup.scala 33:37]
  wire [4:0] _T_1208 = _T_271 ? 5'h14 : _T_1207; // @[Lookup.scala 33:37]
  wire [4:0] _T_1209 = _T_269 ? 5'h14 : _T_1208; // @[Lookup.scala 33:37]
  wire [4:0] _T_1210 = _T_267 ? 5'h14 : _T_1209; // @[Lookup.scala 33:37]
  wire [4:0] _T_1211 = _T_265 ? 5'h14 : _T_1210; // @[Lookup.scala 33:37]
  wire [4:0] _T_1212 = _T_263 ? 5'h14 : _T_1211; // @[Lookup.scala 33:37]
  wire [4:0] _T_1213 = _T_261 ? 5'h14 : _T_1212; // @[Lookup.scala 33:37]
  wire [4:0] _T_1214 = _T_259 ? 5'h14 : _T_1213; // @[Lookup.scala 33:37]
  wire [4:0] _T_1215 = _T_257 ? 5'h14 : _T_1214; // @[Lookup.scala 33:37]
  wire [4:0] _T_1216 = _T_255 ? 5'h14 : _T_1215; // @[Lookup.scala 33:37]
  wire [4:0] _T_1217 = _T_253 ? 5'h14 : _T_1216; // @[Lookup.scala 33:37]
  wire [4:0] _T_1218 = _T_251 ? 5'h14 : _T_1217; // @[Lookup.scala 33:37]
  wire [4:0] _T_1219 = _T_249 ? 5'h14 : _T_1218; // @[Lookup.scala 33:37]
  wire [4:0] _T_1220 = _T_247 ? 5'h1 : _T_1219; // @[Lookup.scala 33:37]
  wire [4:0] _T_1221 = _T_245 ? 5'hc : _T_1220; // @[Lookup.scala 33:37]
  wire [4:0] _T_1222 = _T_243 ? 5'hc : _T_1221; // @[Lookup.scala 33:37]
  wire [4:0] _T_1223 = _T_241 ? 5'hc : _T_1222; // @[Lookup.scala 33:37]
  wire [4:0] _T_1224 = _T_239 ? 5'hc : _T_1223; // @[Lookup.scala 33:37]
  wire [4:0] _T_1225 = _T_237 ? 5'hc : _T_1224; // @[Lookup.scala 33:37]
  wire [4:0] _T_1226 = _T_235 ? 5'hc : _T_1225; // @[Lookup.scala 33:37]
  wire [4:0] _T_1227 = _T_233 ? 5'h5 : _T_1226; // @[Lookup.scala 33:37]
  wire [4:0] _T_1228 = _T_231 ? 5'h5 : _T_1227; // @[Lookup.scala 33:37]
  wire [4:0] _T_1229 = _T_229 ? 5'h5 : _T_1228; // @[Lookup.scala 33:37]
  wire [4:0] _T_1230 = _T_227 ? 5'h5 : _T_1229; // @[Lookup.scala 33:37]
  wire [4:0] _T_1231 = _T_225 ? 5'h5 : _T_1230; // @[Lookup.scala 33:37]
  wire [4:0] _T_1232 = _T_223 ? 5'h5 : _T_1231; // @[Lookup.scala 33:37]
  wire [4:0] _T_1233 = _T_221 ? 5'h5 : _T_1232; // @[Lookup.scala 33:37]
  wire [4:0] _T_1234 = _T_219 ? 5'h5 : _T_1233; // @[Lookup.scala 33:37]
  wire [4:0] _T_1235 = _T_217 ? 5'h5 : _T_1234; // @[Lookup.scala 33:37]
  wire [4:0] _T_1236 = _T_215 ? 5'hf : _T_1235; // @[Lookup.scala 33:37]
  wire [4:0] _T_1237 = _T_213 ? 5'hf : _T_1236; // @[Lookup.scala 33:37]
  wire [4:0] _T_1238 = _T_211 ? 5'h4 : _T_1237; // @[Lookup.scala 33:37]
  wire [4:0] _T_1239 = _T_209 ? 5'h4 : _T_1238; // @[Lookup.scala 33:37]
  wire [4:0] _T_1240 = _T_207 ? 5'h5 : _T_1239; // @[Lookup.scala 33:37]
  wire [4:0] _T_1241 = _T_205 ? 5'hc : _T_1240; // @[Lookup.scala 33:37]
  wire [4:0] _T_1242 = _T_203 ? 5'hc : _T_1241; // @[Lookup.scala 33:37]
  wire [4:0] _T_1243 = _T_201 ? 5'h2 : _T_1242; // @[Lookup.scala 33:37]
  wire [4:0] _T_1244 = _T_199 ? 5'hc : _T_1243; // @[Lookup.scala 33:37]
  wire [4:0] _T_1245 = _T_197 ? 5'hc : _T_1244; // @[Lookup.scala 33:37]
  wire [4:0] _T_1246 = _T_195 ? 5'hc : _T_1245; // @[Lookup.scala 33:37]
  wire [4:0] _T_1247 = _T_193 ? 5'h2 : _T_1246; // @[Lookup.scala 33:37]
  wire [4:0] _T_1248 = _T_191 ? 5'h2 : _T_1247; // @[Lookup.scala 33:37]
  wire [4:0] _T_1249 = _T_189 ? 5'h5 : _T_1248; // @[Lookup.scala 33:37]
  wire [4:0] _T_1250 = _T_187 ? 5'h4 : _T_1249; // @[Lookup.scala 33:37]
  wire [4:0] _T_1251 = _T_185 ? 5'h4 : _T_1250; // @[Lookup.scala 33:37]
  wire [4:0] _T_1252 = _T_183 ? 5'h5 : _T_1251; // @[Lookup.scala 33:37]
  wire [4:0] _T_1253 = _T_181 ? 5'h4 : _T_1252; // @[Lookup.scala 33:37]
  wire [4:0] _T_1254 = _T_179 ? 5'h4 : _T_1253; // @[Lookup.scala 33:37]
  wire [4:0] _T_1255 = _T_177 ? 5'h4 : _T_1254; // @[Lookup.scala 33:37]
  wire [4:0] _T_1256 = _T_175 ? 5'h4 : _T_1255; // @[Lookup.scala 33:37]
  wire [4:0] _T_1257 = _T_173 ? 5'h1 : _T_1256; // @[Lookup.scala 33:37]
  wire [4:0] _T_1258 = _T_171 ? 5'h1 : _T_1257; // @[Lookup.scala 33:37]
  wire [4:0] _T_1259 = _T_169 ? 5'h7 : _T_1258; // @[Lookup.scala 33:37]
  wire [4:0] _T_1260 = _T_167 ? 5'h5 : _T_1259; // @[Lookup.scala 33:37]
  wire [4:0] _T_1261 = _T_165 ? 5'h5 : _T_1260; // @[Lookup.scala 33:37]
  wire [4:0] _T_1262 = _T_163 ? 5'h5 : _T_1261; // @[Lookup.scala 33:37]
  wire [4:0] _T_1263 = _T_161 ? 5'h5 : _T_1262; // @[Lookup.scala 33:37]
  wire [4:0] _T_1264 = _T_159 ? 5'h5 : _T_1263; // @[Lookup.scala 33:37]
  wire [4:0] _T_1265 = _T_157 ? 5'h5 : _T_1264; // @[Lookup.scala 33:37]
  wire [4:0] _T_1266 = _T_155 ? 5'h4 : _T_1265; // @[Lookup.scala 33:37]
  wire [4:0] _T_1267 = _T_153 ? 5'h4 : _T_1266; // @[Lookup.scala 33:37]
  wire [4:0] _T_1268 = _T_151 ? 5'h4 : _T_1267; // @[Lookup.scala 33:37]
  wire [4:0] _T_1269 = _T_149 ? 5'h4 : _T_1268; // @[Lookup.scala 33:37]
  wire [4:0] _T_1270 = _T_147 ? 5'h4 : _T_1269; // @[Lookup.scala 33:37]
  wire [4:0] _T_1271 = _T_145 ? 5'h4 : _T_1270; // @[Lookup.scala 33:37]
  wire [4:0] _T_1272 = _T_143 ? 5'h4 : _T_1271; // @[Lookup.scala 33:37]
  wire [4:0] _T_1273 = _T_141 ? 5'h4 : _T_1272; // @[Lookup.scala 33:37]
  wire [4:0] _T_1274 = _T_139 ? 5'h4 : _T_1273; // @[Lookup.scala 33:37]
  wire [4:0] _T_1275 = _T_137 ? 5'h2 : _T_1274; // @[Lookup.scala 33:37]
  wire [4:0] _T_1276 = _T_135 ? 5'h2 : _T_1275; // @[Lookup.scala 33:37]
  wire [4:0] _T_1277 = _T_133 ? 5'h4 : _T_1276; // @[Lookup.scala 33:37]
  wire [4:0] _T_1278 = _T_131 ? 5'h4 : _T_1277; // @[Lookup.scala 33:37]
  wire [4:0] _T_1279 = _T_129 ? 5'h4 : _T_1278; // @[Lookup.scala 33:37]
  wire [4:0] _T_1280 = _T_127 ? 5'h0 : _T_1279; // @[Lookup.scala 33:37]
  wire [4:0] _T_1281 = _T_125 ? 5'h5 : _T_1280; // @[Lookup.scala 33:37]
  wire [4:0] _T_1282 = _T_123 ? 5'h5 : _T_1281; // @[Lookup.scala 33:37]
  wire [4:0] _T_1283 = _T_121 ? 5'h5 : _T_1282; // @[Lookup.scala 33:37]
  wire [4:0] _T_1284 = _T_119 ? 5'h5 : _T_1283; // @[Lookup.scala 33:37]
  wire [4:0] _T_1285 = _T_117 ? 5'h5 : _T_1284; // @[Lookup.scala 33:37]
  wire [4:0] _T_1286 = _T_115 ? 5'h5 : _T_1285; // @[Lookup.scala 33:37]
  wire [4:0] _T_1287 = _T_113 ? 5'h5 : _T_1286; // @[Lookup.scala 33:37]
  wire [4:0] _T_1288 = _T_111 ? 5'h5 : _T_1287; // @[Lookup.scala 33:37]
  wire [4:0] _T_1289 = _T_109 ? 5'h5 : _T_1288; // @[Lookup.scala 33:37]
  wire [4:0] _T_1290 = _T_107 ? 5'h5 : _T_1289; // @[Lookup.scala 33:37]
  wire [4:0] _T_1291 = _T_105 ? 5'h5 : _T_1290; // @[Lookup.scala 33:37]
  wire [4:0] _T_1292 = _T_103 ? 5'h5 : _T_1291; // @[Lookup.scala 33:37]
  wire [4:0] _T_1293 = _T_101 ? 5'h5 : _T_1292; // @[Lookup.scala 33:37]
  wire [4:0] _T_1294 = _T_99 ? 5'h4 : _T_1293; // @[Lookup.scala 33:37]
  wire [4:0] _T_1295 = _T_97 ? 5'h2 : _T_1294; // @[Lookup.scala 33:37]
  wire [4:0] _T_1296 = _T_95 ? 5'h4 : _T_1295; // @[Lookup.scala 33:37]
  wire [4:0] _T_1297 = _T_93 ? 5'h4 : _T_1296; // @[Lookup.scala 33:37]
  wire [4:0] _T_1298 = _T_91 ? 5'h5 : _T_1297; // @[Lookup.scala 33:37]
  wire [4:0] _T_1299 = _T_89 ? 5'h5 : _T_1298; // @[Lookup.scala 33:37]
  wire [4:0] _T_1300 = _T_87 ? 5'h5 : _T_1299; // @[Lookup.scala 33:37]
  wire [4:0] _T_1301 = _T_85 ? 5'h5 : _T_1300; // @[Lookup.scala 33:37]
  wire [4:0] _T_1302 = _T_83 ? 5'h5 : _T_1301; // @[Lookup.scala 33:37]
  wire [4:0] _T_1303 = _T_81 ? 5'h4 : _T_1302; // @[Lookup.scala 33:37]
  wire [4:0] _T_1304 = _T_79 ? 5'h4 : _T_1303; // @[Lookup.scala 33:37]
  wire [4:0] _T_1305 = _T_77 ? 5'h4 : _T_1304; // @[Lookup.scala 33:37]
  wire [4:0] _T_1306 = _T_75 ? 5'h4 : _T_1305; // @[Lookup.scala 33:37]
  wire [4:0] _T_1307 = _T_73 ? 5'h2 : _T_1306; // @[Lookup.scala 33:37]
  wire [4:0] _T_1308 = _T_71 ? 5'h2 : _T_1307; // @[Lookup.scala 33:37]
  wire [4:0] _T_1309 = _T_69 ? 5'h2 : _T_1308; // @[Lookup.scala 33:37]
  wire [4:0] _T_1310 = _T_67 ? 5'h4 : _T_1309; // @[Lookup.scala 33:37]
  wire [4:0] _T_1311 = _T_65 ? 5'h4 : _T_1310; // @[Lookup.scala 33:37]
  wire [4:0] _T_1312 = _T_63 ? 5'h4 : _T_1311; // @[Lookup.scala 33:37]
  wire [4:0] _T_1313 = _T_61 ? 5'h4 : _T_1312; // @[Lookup.scala 33:37]
  wire [4:0] _T_1314 = _T_59 ? 5'h4 : _T_1313; // @[Lookup.scala 33:37]
  wire [4:0] _T_1315 = _T_57 ? 5'h1 : _T_1314; // @[Lookup.scala 33:37]
  wire [4:0] _T_1316 = _T_55 ? 5'h1 : _T_1315; // @[Lookup.scala 33:37]
  wire [4:0] _T_1317 = _T_53 ? 5'h1 : _T_1316; // @[Lookup.scala 33:37]
  wire [4:0] _T_1318 = _T_51 ? 5'h1 : _T_1317; // @[Lookup.scala 33:37]
  wire [4:0] _T_1319 = _T_49 ? 5'h1 : _T_1318; // @[Lookup.scala 33:37]
  wire [4:0] _T_1320 = _T_47 ? 5'h1 : _T_1319; // @[Lookup.scala 33:37]
  wire [4:0] _T_1321 = _T_45 ? 5'h4 : _T_1320; // @[Lookup.scala 33:37]
  wire [4:0] _T_1322 = _T_43 ? 5'h7 : _T_1321; // @[Lookup.scala 33:37]
  wire [4:0] _T_1323 = _T_41 ? 5'h6 : _T_1322; // @[Lookup.scala 33:37]
  wire [4:0] _T_1324 = _T_39 ? 5'h6 : _T_1323; // @[Lookup.scala 33:37]
  wire [4:0] _T_1325 = _T_37 ? 5'h5 : _T_1324; // @[Lookup.scala 33:37]
  wire [4:0] _T_1326 = _T_35 ? 5'h5 : _T_1325; // @[Lookup.scala 33:37]
  wire [4:0] _T_1327 = _T_33 ? 5'h5 : _T_1326; // @[Lookup.scala 33:37]
  wire [4:0] _T_1328 = _T_31 ? 5'h5 : _T_1327; // @[Lookup.scala 33:37]
  wire [4:0] _T_1329 = _T_29 ? 5'h5 : _T_1328; // @[Lookup.scala 33:37]
  wire [4:0] _T_1330 = _T_27 ? 5'h5 : _T_1329; // @[Lookup.scala 33:37]
  wire [4:0] _T_1331 = _T_25 ? 5'h5 : _T_1330; // @[Lookup.scala 33:37]
  wire [4:0] _T_1332 = _T_23 ? 5'h5 : _T_1331; // @[Lookup.scala 33:37]
  wire [4:0] _T_1333 = _T_21 ? 5'h5 : _T_1332; // @[Lookup.scala 33:37]
  wire [4:0] _T_1334 = _T_19 ? 5'h5 : _T_1333; // @[Lookup.scala 33:37]
  wire [4:0] _T_1335 = _T_17 ? 5'h4 : _T_1334; // @[Lookup.scala 33:37]
  wire [4:0] _T_1336 = _T_15 ? 5'h4 : _T_1335; // @[Lookup.scala 33:37]
  wire [4:0] _T_1337 = _T_13 ? 5'h4 : _T_1336; // @[Lookup.scala 33:37]
  wire [4:0] _T_1338 = _T_11 ? 5'h4 : _T_1337; // @[Lookup.scala 33:37]
  wire [4:0] _T_1339 = _T_9 ? 5'h4 : _T_1338; // @[Lookup.scala 33:37]
  wire [4:0] _T_1340 = _T_7 ? 5'h4 : _T_1339; // @[Lookup.scala 33:37]
  wire [4:0] _T_1341 = _T_5 ? 5'h4 : _T_1340; // @[Lookup.scala 33:37]
  wire [4:0] _T_1342 = _T_3 ? 5'h4 : _T_1341; // @[Lookup.scala 33:37]
  wire [4:0] decodeList_0 = _T_1 ? 5'h4 : _T_1342; // @[Lookup.scala 33:37]
  wire [3:0] _T_1343 = _T_895 ? 4'h2 : 4'h1; // @[Lookup.scala 33:37]
  wire [3:0] _T_1344 = _T_893 ? 4'h2 : _T_1343; // @[Lookup.scala 33:37]
  wire [3:0] _T_1345 = _T_891 ? 4'h2 : _T_1344; // @[Lookup.scala 33:37]
  wire [3:0] _T_1346 = _T_889 ? 4'h2 : _T_1345; // @[Lookup.scala 33:37]
  wire [3:0] _T_1347 = _T_887 ? 4'h2 : _T_1346; // @[Lookup.scala 33:37]
  wire [3:0] _T_1348 = _T_885 ? 4'h2 : _T_1347; // @[Lookup.scala 33:37]
  wire [3:0] _T_1349 = _T_883 ? 4'h2 : _T_1348; // @[Lookup.scala 33:37]
  wire [3:0] _T_1350 = _T_881 ? 4'h2 : _T_1349; // @[Lookup.scala 33:37]
  wire [3:0] _T_1351 = _T_879 ? 4'h2 : _T_1350; // @[Lookup.scala 33:37]
  wire [3:0] _T_1352 = _T_877 ? 4'h2 : _T_1351; // @[Lookup.scala 33:37]
  wire [3:0] _T_1353 = _T_875 ? 4'h2 : _T_1352; // @[Lookup.scala 33:37]
  wire [3:0] _T_1354 = _T_873 ? 4'h2 : _T_1353; // @[Lookup.scala 33:37]
  wire [3:0] _T_1355 = _T_871 ? 4'h2 : _T_1354; // @[Lookup.scala 33:37]
  wire [3:0] _T_1356 = _T_869 ? 4'h2 : _T_1355; // @[Lookup.scala 33:37]
  wire [3:0] _T_1357 = _T_867 ? 4'h2 : _T_1356; // @[Lookup.scala 33:37]
  wire [3:0] _T_1358 = _T_865 ? 4'h2 : _T_1357; // @[Lookup.scala 33:37]
  wire [3:0] _T_1359 = _T_863 ? 4'h2 : _T_1358; // @[Lookup.scala 33:37]
  wire [3:0] _T_1360 = _T_861 ? 4'h2 : _T_1359; // @[Lookup.scala 33:37]
  wire [3:0] _T_1361 = _T_859 ? 4'h2 : _T_1360; // @[Lookup.scala 33:37]
  wire [3:0] _T_1362 = _T_857 ? 4'h2 : _T_1361; // @[Lookup.scala 33:37]
  wire [3:0] _T_1363 = _T_855 ? 4'h2 : _T_1362; // @[Lookup.scala 33:37]
  wire [3:0] _T_1364 = _T_853 ? 4'h2 : _T_1363; // @[Lookup.scala 33:37]
  wire [3:0] _T_1365 = _T_851 ? 4'h2 : _T_1364; // @[Lookup.scala 33:37]
  wire [3:0] _T_1366 = _T_849 ? 4'h2 : _T_1365; // @[Lookup.scala 33:37]
  wire [3:0] _T_1367 = _T_847 ? 4'h2 : _T_1366; // @[Lookup.scala 33:37]
  wire [3:0] _T_1368 = _T_845 ? 4'h2 : _T_1367; // @[Lookup.scala 33:37]
  wire [3:0] _T_1369 = _T_843 ? 4'h2 : _T_1368; // @[Lookup.scala 33:37]
  wire [3:0] _T_1370 = _T_841 ? 4'h2 : _T_1369; // @[Lookup.scala 33:37]
  wire [3:0] _T_1371 = _T_839 ? 4'h2 : _T_1370; // @[Lookup.scala 33:37]
  wire [3:0] _T_1372 = _T_837 ? 4'h2 : _T_1371; // @[Lookup.scala 33:37]
  wire [3:0] _T_1373 = _T_835 ? 4'h2 : _T_1372; // @[Lookup.scala 33:37]
  wire [3:0] _T_1374 = _T_833 ? 4'h2 : _T_1373; // @[Lookup.scala 33:37]
  wire [3:0] _T_1375 = _T_831 ? 4'h2 : _T_1374; // @[Lookup.scala 33:37]
  wire [3:0] _T_1376 = _T_829 ? 4'h2 : _T_1375; // @[Lookup.scala 33:37]
  wire [3:0] _T_1377 = _T_827 ? 4'h2 : _T_1376; // @[Lookup.scala 33:37]
  wire [3:0] _T_1378 = _T_825 ? 4'h2 : _T_1377; // @[Lookup.scala 33:37]
  wire [3:0] _T_1379 = _T_823 ? 4'h2 : _T_1378; // @[Lookup.scala 33:37]
  wire [3:0] _T_1380 = _T_821 ? 4'h2 : _T_1379; // @[Lookup.scala 33:37]
  wire [3:0] _T_1381 = _T_819 ? 4'h2 : _T_1380; // @[Lookup.scala 33:37]
  wire [3:0] _T_1382 = _T_817 ? 4'h2 : _T_1381; // @[Lookup.scala 33:37]
  wire [3:0] _T_1383 = _T_815 ? 4'h2 : _T_1382; // @[Lookup.scala 33:37]
  wire [3:0] _T_1384 = _T_813 ? 4'h2 : _T_1383; // @[Lookup.scala 33:37]
  wire [3:0] _T_1385 = _T_811 ? 4'h2 : _T_1384; // @[Lookup.scala 33:37]
  wire [3:0] _T_1386 = _T_809 ? 4'h2 : _T_1385; // @[Lookup.scala 33:37]
  wire [3:0] _T_1387 = _T_807 ? 4'h2 : _T_1386; // @[Lookup.scala 33:37]
  wire [3:0] _T_1388 = _T_805 ? 4'h2 : _T_1387; // @[Lookup.scala 33:37]
  wire [3:0] _T_1389 = _T_803 ? 4'h2 : _T_1388; // @[Lookup.scala 33:37]
  wire [3:0] _T_1390 = _T_801 ? 4'h2 : _T_1389; // @[Lookup.scala 33:37]
  wire [3:0] _T_1391 = _T_799 ? 4'h2 : _T_1390; // @[Lookup.scala 33:37]
  wire [3:0] _T_1392 = _T_797 ? 4'h2 : _T_1391; // @[Lookup.scala 33:37]
  wire [3:0] _T_1393 = _T_795 ? 4'h2 : _T_1392; // @[Lookup.scala 33:37]
  wire [3:0] _T_1394 = _T_793 ? 4'h2 : _T_1393; // @[Lookup.scala 33:37]
  wire [3:0] _T_1395 = _T_791 ? 4'h2 : _T_1394; // @[Lookup.scala 33:37]
  wire [3:0] _T_1396 = _T_789 ? 4'h2 : _T_1395; // @[Lookup.scala 33:37]
  wire [3:0] _T_1397 = _T_787 ? 4'h2 : _T_1396; // @[Lookup.scala 33:37]
  wire [3:0] _T_1398 = _T_785 ? 4'h2 : _T_1397; // @[Lookup.scala 33:37]
  wire [3:0] _T_1399 = _T_783 ? 4'h2 : _T_1398; // @[Lookup.scala 33:37]
  wire [3:0] _T_1400 = _T_781 ? 4'h2 : _T_1399; // @[Lookup.scala 33:37]
  wire [3:0] _T_1401 = _T_779 ? 4'h2 : _T_1400; // @[Lookup.scala 33:37]
  wire [3:0] _T_1402 = _T_777 ? 4'h2 : _T_1401; // @[Lookup.scala 33:37]
  wire [3:0] _T_1403 = _T_775 ? 4'h2 : _T_1402; // @[Lookup.scala 33:37]
  wire [3:0] _T_1404 = _T_773 ? 4'h2 : _T_1403; // @[Lookup.scala 33:37]
  wire [3:0] _T_1405 = _T_771 ? 4'h2 : _T_1404; // @[Lookup.scala 33:37]
  wire [3:0] _T_1406 = _T_769 ? 4'h2 : _T_1405; // @[Lookup.scala 33:37]
  wire [3:0] _T_1407 = _T_767 ? 4'h2 : _T_1406; // @[Lookup.scala 33:37]
  wire [3:0] _T_1408 = _T_765 ? 4'h2 : _T_1407; // @[Lookup.scala 33:37]
  wire [3:0] _T_1409 = _T_763 ? 4'h2 : _T_1408; // @[Lookup.scala 33:37]
  wire [3:0] _T_1410 = _T_761 ? 4'h2 : _T_1409; // @[Lookup.scala 33:37]
  wire [3:0] _T_1411 = _T_759 ? 4'h2 : _T_1410; // @[Lookup.scala 33:37]
  wire [3:0] _T_1412 = _T_757 ? 4'h2 : _T_1411; // @[Lookup.scala 33:37]
  wire [3:0] _T_1413 = _T_755 ? 4'h2 : _T_1412; // @[Lookup.scala 33:37]
  wire [3:0] _T_1414 = _T_753 ? 4'h2 : _T_1413; // @[Lookup.scala 33:37]
  wire [3:0] _T_1415 = _T_751 ? 4'h2 : _T_1414; // @[Lookup.scala 33:37]
  wire [3:0] _T_1416 = _T_749 ? 4'h2 : _T_1415; // @[Lookup.scala 33:37]
  wire [3:0] _T_1417 = _T_747 ? 4'h2 : _T_1416; // @[Lookup.scala 33:37]
  wire [3:0] _T_1418 = _T_745 ? 4'h2 : _T_1417; // @[Lookup.scala 33:37]
  wire [3:0] _T_1419 = _T_743 ? 4'h2 : _T_1418; // @[Lookup.scala 33:37]
  wire [3:0] _T_1420 = _T_741 ? 4'h2 : _T_1419; // @[Lookup.scala 33:37]
  wire [3:0] _T_1421 = _T_739 ? 4'h2 : _T_1420; // @[Lookup.scala 33:37]
  wire [3:0] _T_1422 = _T_737 ? 4'h2 : _T_1421; // @[Lookup.scala 33:37]
  wire [3:0] _T_1423 = _T_735 ? 4'h2 : _T_1422; // @[Lookup.scala 33:37]
  wire [3:0] _T_1424 = _T_733 ? 4'h2 : _T_1423; // @[Lookup.scala 33:37]
  wire [3:0] _T_1425 = _T_731 ? 4'h2 : _T_1424; // @[Lookup.scala 33:37]
  wire [3:0] _T_1426 = _T_729 ? 4'h2 : _T_1425; // @[Lookup.scala 33:37]
  wire [3:0] _T_1427 = _T_727 ? 4'h2 : _T_1426; // @[Lookup.scala 33:37]
  wire [3:0] _T_1428 = _T_725 ? 4'h2 : _T_1427; // @[Lookup.scala 33:37]
  wire [3:0] _T_1429 = _T_723 ? 4'h2 : _T_1428; // @[Lookup.scala 33:37]
  wire [3:0] _T_1430 = _T_721 ? 4'h2 : _T_1429; // @[Lookup.scala 33:37]
  wire [3:0] _T_1431 = _T_719 ? 4'h2 : _T_1430; // @[Lookup.scala 33:37]
  wire [3:0] _T_1432 = _T_717 ? 4'h2 : _T_1431; // @[Lookup.scala 33:37]
  wire [3:0] _T_1433 = _T_715 ? 4'h2 : _T_1432; // @[Lookup.scala 33:37]
  wire [3:0] _T_1434 = _T_713 ? 4'h2 : _T_1433; // @[Lookup.scala 33:37]
  wire [3:0] _T_1435 = _T_711 ? 4'h2 : _T_1434; // @[Lookup.scala 33:37]
  wire [3:0] _T_1436 = _T_709 ? 4'h2 : _T_1435; // @[Lookup.scala 33:37]
  wire [3:0] _T_1437 = _T_707 ? 4'h2 : _T_1436; // @[Lookup.scala 33:37]
  wire [3:0] _T_1438 = _T_705 ? 4'h2 : _T_1437; // @[Lookup.scala 33:37]
  wire [3:0] _T_1439 = _T_703 ? 4'h2 : _T_1438; // @[Lookup.scala 33:37]
  wire [3:0] _T_1440 = _T_701 ? 4'h2 : _T_1439; // @[Lookup.scala 33:37]
  wire [3:0] _T_1441 = _T_699 ? 4'h2 : _T_1440; // @[Lookup.scala 33:37]
  wire [3:0] _T_1442 = _T_697 ? 4'h2 : _T_1441; // @[Lookup.scala 33:37]
  wire [3:0] _T_1443 = _T_695 ? 4'h2 : _T_1442; // @[Lookup.scala 33:37]
  wire [3:0] _T_1444 = _T_693 ? 4'h2 : _T_1443; // @[Lookup.scala 33:37]
  wire [3:0] _T_1445 = _T_691 ? 4'h2 : _T_1444; // @[Lookup.scala 33:37]
  wire [3:0] _T_1446 = _T_689 ? 4'h2 : _T_1445; // @[Lookup.scala 33:37]
  wire [3:0] _T_1447 = _T_687 ? 4'h2 : _T_1446; // @[Lookup.scala 33:37]
  wire [3:0] _T_1448 = _T_685 ? 4'h2 : _T_1447; // @[Lookup.scala 33:37]
  wire [3:0] _T_1449 = _T_683 ? 4'h2 : _T_1448; // @[Lookup.scala 33:37]
  wire [3:0] _T_1450 = _T_681 ? 4'h2 : _T_1449; // @[Lookup.scala 33:37]
  wire [3:0] _T_1451 = _T_679 ? 4'h2 : _T_1450; // @[Lookup.scala 33:37]
  wire [3:0] _T_1452 = _T_677 ? 4'h2 : _T_1451; // @[Lookup.scala 33:37]
  wire [3:0] _T_1453 = _T_675 ? 4'h2 : _T_1452; // @[Lookup.scala 33:37]
  wire [3:0] _T_1454 = _T_673 ? 4'h2 : _T_1453; // @[Lookup.scala 33:37]
  wire [3:0] _T_1455 = _T_671 ? 4'h2 : _T_1454; // @[Lookup.scala 33:37]
  wire [3:0] _T_1456 = _T_669 ? 4'h2 : _T_1455; // @[Lookup.scala 33:37]
  wire [3:0] _T_1457 = _T_667 ? 4'h2 : _T_1456; // @[Lookup.scala 33:37]
  wire [3:0] _T_1458 = _T_665 ? 4'h2 : _T_1457; // @[Lookup.scala 33:37]
  wire [3:0] _T_1459 = _T_663 ? 4'h2 : _T_1458; // @[Lookup.scala 33:37]
  wire [3:0] _T_1460 = _T_661 ? 4'h2 : _T_1459; // @[Lookup.scala 33:37]
  wire [3:0] _T_1461 = _T_659 ? 4'h2 : _T_1460; // @[Lookup.scala 33:37]
  wire [3:0] _T_1462 = _T_657 ? 4'h2 : _T_1461; // @[Lookup.scala 33:37]
  wire [3:0] _T_1463 = _T_655 ? 4'h2 : _T_1462; // @[Lookup.scala 33:37]
  wire [3:0] _T_1464 = _T_653 ? 4'h2 : _T_1463; // @[Lookup.scala 33:37]
  wire [3:0] _T_1465 = _T_651 ? 4'h2 : _T_1464; // @[Lookup.scala 33:37]
  wire [3:0] _T_1466 = _T_649 ? 4'h2 : _T_1465; // @[Lookup.scala 33:37]
  wire [3:0] _T_1467 = _T_647 ? 4'h2 : _T_1466; // @[Lookup.scala 33:37]
  wire [3:0] _T_1468 = _T_645 ? 4'h2 : _T_1467; // @[Lookup.scala 33:37]
  wire [3:0] _T_1469 = _T_643 ? 4'h2 : _T_1468; // @[Lookup.scala 33:37]
  wire [3:0] _T_1470 = _T_641 ? 4'h2 : _T_1469; // @[Lookup.scala 33:37]
  wire [3:0] _T_1471 = _T_639 ? 4'h2 : _T_1470; // @[Lookup.scala 33:37]
  wire [3:0] _T_1472 = _T_637 ? 4'h2 : _T_1471; // @[Lookup.scala 33:37]
  wire [3:0] _T_1473 = _T_635 ? 4'h2 : _T_1472; // @[Lookup.scala 33:37]
  wire [3:0] _T_1474 = _T_633 ? 4'h2 : _T_1473; // @[Lookup.scala 33:37]
  wire [3:0] _T_1475 = _T_631 ? 4'h2 : _T_1474; // @[Lookup.scala 33:37]
  wire [3:0] _T_1476 = _T_629 ? 4'h2 : _T_1475; // @[Lookup.scala 33:37]
  wire [3:0] _T_1477 = _T_627 ? 4'h2 : _T_1476; // @[Lookup.scala 33:37]
  wire [3:0] _T_1478 = _T_625 ? 4'h2 : _T_1477; // @[Lookup.scala 33:37]
  wire [3:0] _T_1479 = _T_623 ? 4'h2 : _T_1478; // @[Lookup.scala 33:37]
  wire [3:0] _T_1480 = _T_621 ? 4'h2 : _T_1479; // @[Lookup.scala 33:37]
  wire [3:0] _T_1481 = _T_619 ? 4'h2 : _T_1480; // @[Lookup.scala 33:37]
  wire [3:0] _T_1482 = _T_617 ? 4'h2 : _T_1481; // @[Lookup.scala 33:37]
  wire [3:0] _T_1483 = _T_615 ? 4'h2 : _T_1482; // @[Lookup.scala 33:37]
  wire [3:0] _T_1484 = _T_613 ? 4'h2 : _T_1483; // @[Lookup.scala 33:37]
  wire [3:0] _T_1485 = _T_611 ? 4'h2 : _T_1484; // @[Lookup.scala 33:37]
  wire [3:0] _T_1486 = _T_609 ? 4'h2 : _T_1485; // @[Lookup.scala 33:37]
  wire [3:0] _T_1487 = _T_607 ? 4'h2 : _T_1486; // @[Lookup.scala 33:37]
  wire [3:0] _T_1488 = _T_605 ? 4'h2 : _T_1487; // @[Lookup.scala 33:37]
  wire [3:0] _T_1489 = _T_603 ? 4'h2 : _T_1488; // @[Lookup.scala 33:37]
  wire [3:0] _T_1490 = _T_601 ? 4'h2 : _T_1489; // @[Lookup.scala 33:37]
  wire [3:0] _T_1491 = _T_599 ? 4'h2 : _T_1490; // @[Lookup.scala 33:37]
  wire [3:0] _T_1492 = _T_597 ? 4'h2 : _T_1491; // @[Lookup.scala 33:37]
  wire [3:0] _T_1493 = _T_595 ? 4'h2 : _T_1492; // @[Lookup.scala 33:37]
  wire [3:0] _T_1494 = _T_593 ? 4'h2 : _T_1493; // @[Lookup.scala 33:37]
  wire [3:0] _T_1495 = _T_591 ? 4'h2 : _T_1494; // @[Lookup.scala 33:37]
  wire [3:0] _T_1496 = _T_589 ? 4'h2 : _T_1495; // @[Lookup.scala 33:37]
  wire [3:0] _T_1497 = _T_587 ? 4'h2 : _T_1496; // @[Lookup.scala 33:37]
  wire [3:0] _T_1498 = _T_585 ? 4'h2 : _T_1497; // @[Lookup.scala 33:37]
  wire [3:0] _T_1499 = _T_583 ? 4'h2 : _T_1498; // @[Lookup.scala 33:37]
  wire [3:0] _T_1500 = _T_581 ? 4'h2 : _T_1499; // @[Lookup.scala 33:37]
  wire [3:0] _T_1501 = _T_579 ? 4'h2 : _T_1500; // @[Lookup.scala 33:37]
  wire [3:0] _T_1502 = _T_577 ? 4'h2 : _T_1501; // @[Lookup.scala 33:37]
  wire [3:0] _T_1503 = _T_575 ? 4'h2 : _T_1502; // @[Lookup.scala 33:37]
  wire [3:0] _T_1504 = _T_573 ? 4'h2 : _T_1503; // @[Lookup.scala 33:37]
  wire [3:0] _T_1505 = _T_571 ? 4'h2 : _T_1504; // @[Lookup.scala 33:37]
  wire [3:0] _T_1506 = _T_569 ? 4'h2 : _T_1505; // @[Lookup.scala 33:37]
  wire [3:0] _T_1507 = _T_567 ? 4'h2 : _T_1506; // @[Lookup.scala 33:37]
  wire [3:0] _T_1508 = _T_565 ? 4'h2 : _T_1507; // @[Lookup.scala 33:37]
  wire [3:0] _T_1509 = _T_563 ? 4'h2 : _T_1508; // @[Lookup.scala 33:37]
  wire [3:0] _T_1510 = _T_561 ? 4'h2 : _T_1509; // @[Lookup.scala 33:37]
  wire [3:0] _T_1511 = _T_559 ? 4'h2 : _T_1510; // @[Lookup.scala 33:37]
  wire [3:0] _T_1512 = _T_557 ? 4'h2 : _T_1511; // @[Lookup.scala 33:37]
  wire [3:0] _T_1513 = _T_555 ? 4'h2 : _T_1512; // @[Lookup.scala 33:37]
  wire [3:0] _T_1514 = _T_553 ? 4'h2 : _T_1513; // @[Lookup.scala 33:37]
  wire [3:0] _T_1515 = _T_551 ? 4'h2 : _T_1514; // @[Lookup.scala 33:37]
  wire [3:0] _T_1516 = _T_549 ? 4'h2 : _T_1515; // @[Lookup.scala 33:37]
  wire [3:0] _T_1517 = _T_547 ? 4'h2 : _T_1516; // @[Lookup.scala 33:37]
  wire [3:0] _T_1518 = _T_545 ? 4'h2 : _T_1517; // @[Lookup.scala 33:37]
  wire [3:0] _T_1519 = _T_543 ? 4'h2 : _T_1518; // @[Lookup.scala 33:37]
  wire [3:0] _T_1520 = _T_541 ? 4'h2 : _T_1519; // @[Lookup.scala 33:37]
  wire [3:0] _T_1521 = _T_539 ? 4'h2 : _T_1520; // @[Lookup.scala 33:37]
  wire [3:0] _T_1522 = _T_537 ? 4'h2 : _T_1521; // @[Lookup.scala 33:37]
  wire [3:0] _T_1523 = _T_535 ? 4'h2 : _T_1522; // @[Lookup.scala 33:37]
  wire [3:0] _T_1524 = _T_533 ? 4'h2 : _T_1523; // @[Lookup.scala 33:37]
  wire [3:0] _T_1525 = _T_531 ? 4'h2 : _T_1524; // @[Lookup.scala 33:37]
  wire [3:0] _T_1526 = _T_529 ? 4'h2 : _T_1525; // @[Lookup.scala 33:37]
  wire [3:0] _T_1527 = _T_527 ? 4'h2 : _T_1526; // @[Lookup.scala 33:37]
  wire [3:0] _T_1528 = _T_525 ? 4'h2 : _T_1527; // @[Lookup.scala 33:37]
  wire [3:0] _T_1529 = _T_523 ? 4'h2 : _T_1528; // @[Lookup.scala 33:37]
  wire [3:0] _T_1530 = _T_521 ? 4'h2 : _T_1529; // @[Lookup.scala 33:37]
  wire [3:0] _T_1531 = _T_519 ? 4'h2 : _T_1530; // @[Lookup.scala 33:37]
  wire [3:0] _T_1532 = _T_517 ? 4'h2 : _T_1531; // @[Lookup.scala 33:37]
  wire [3:0] _T_1533 = _T_515 ? 4'h2 : _T_1532; // @[Lookup.scala 33:37]
  wire [3:0] _T_1534 = _T_513 ? 4'h2 : _T_1533; // @[Lookup.scala 33:37]
  wire [3:0] _T_1535 = _T_511 ? 4'h2 : _T_1534; // @[Lookup.scala 33:37]
  wire [3:0] _T_1536 = _T_509 ? 4'h2 : _T_1535; // @[Lookup.scala 33:37]
  wire [3:0] _T_1537 = _T_507 ? 4'h2 : _T_1536; // @[Lookup.scala 33:37]
  wire [3:0] _T_1538 = _T_505 ? 4'h2 : _T_1537; // @[Lookup.scala 33:37]
  wire [3:0] _T_1539 = _T_503 ? 4'h2 : _T_1538; // @[Lookup.scala 33:37]
  wire [3:0] _T_1540 = _T_501 ? 4'h2 : _T_1539; // @[Lookup.scala 33:37]
  wire [3:0] _T_1541 = _T_499 ? 4'h2 : _T_1540; // @[Lookup.scala 33:37]
  wire [3:0] _T_1542 = _T_497 ? 4'h2 : _T_1541; // @[Lookup.scala 33:37]
  wire [3:0] _T_1543 = _T_495 ? 4'h2 : _T_1542; // @[Lookup.scala 33:37]
  wire [3:0] _T_1544 = _T_493 ? 4'h2 : _T_1543; // @[Lookup.scala 33:37]
  wire [3:0] _T_1545 = _T_491 ? 4'h2 : _T_1544; // @[Lookup.scala 33:37]
  wire [3:0] _T_1546 = _T_489 ? 4'h2 : _T_1545; // @[Lookup.scala 33:37]
  wire [3:0] _T_1547 = _T_487 ? 4'h2 : _T_1546; // @[Lookup.scala 33:37]
  wire [3:0] _T_1548 = _T_485 ? 4'h2 : _T_1547; // @[Lookup.scala 33:37]
  wire [3:0] _T_1549 = _T_483 ? 4'h2 : _T_1548; // @[Lookup.scala 33:37]
  wire [3:0] _T_1550 = _T_481 ? 4'h2 : _T_1549; // @[Lookup.scala 33:37]
  wire [3:0] _T_1551 = _T_479 ? 4'h2 : _T_1550; // @[Lookup.scala 33:37]
  wire [3:0] _T_1552 = _T_477 ? 4'h2 : _T_1551; // @[Lookup.scala 33:37]
  wire [3:0] _T_1553 = _T_475 ? 4'h2 : _T_1552; // @[Lookup.scala 33:37]
  wire [3:0] _T_1554 = _T_473 ? 4'h2 : _T_1553; // @[Lookup.scala 33:37]
  wire [3:0] _T_1555 = _T_471 ? 4'h2 : _T_1554; // @[Lookup.scala 33:37]
  wire [3:0] _T_1556 = _T_469 ? 4'h2 : _T_1555; // @[Lookup.scala 33:37]
  wire [3:0] _T_1557 = _T_467 ? 4'h2 : _T_1556; // @[Lookup.scala 33:37]
  wire [3:0] _T_1558 = _T_465 ? 4'h2 : _T_1557; // @[Lookup.scala 33:37]
  wire [3:0] _T_1559 = _T_463 ? 4'h2 : _T_1558; // @[Lookup.scala 33:37]
  wire [3:0] _T_1560 = _T_461 ? 4'h2 : _T_1559; // @[Lookup.scala 33:37]
  wire [3:0] _T_1561 = _T_459 ? 4'h2 : _T_1560; // @[Lookup.scala 33:37]
  wire [3:0] _T_1562 = _T_457 ? 4'h2 : _T_1561; // @[Lookup.scala 33:37]
  wire [3:0] _T_1563 = _T_455 ? 4'h2 : _T_1562; // @[Lookup.scala 33:37]
  wire [3:0] _T_1564 = _T_453 ? 4'h2 : _T_1563; // @[Lookup.scala 33:37]
  wire [3:0] _T_1565 = _T_451 ? 4'h2 : _T_1564; // @[Lookup.scala 33:37]
  wire [3:0] _T_1566 = _T_449 ? 4'h2 : _T_1565; // @[Lookup.scala 33:37]
  wire [3:0] _T_1567 = _T_447 ? 4'h2 : _T_1566; // @[Lookup.scala 33:37]
  wire [3:0] _T_1568 = _T_445 ? 4'h2 : _T_1567; // @[Lookup.scala 33:37]
  wire [3:0] _T_1569 = _T_443 ? 4'h2 : _T_1568; // @[Lookup.scala 33:37]
  wire [3:0] _T_1570 = _T_441 ? 4'h2 : _T_1569; // @[Lookup.scala 33:37]
  wire [3:0] _T_1571 = _T_439 ? 4'h2 : _T_1570; // @[Lookup.scala 33:37]
  wire [3:0] _T_1572 = _T_437 ? 4'h2 : _T_1571; // @[Lookup.scala 33:37]
  wire [3:0] _T_1573 = _T_435 ? 4'h2 : _T_1572; // @[Lookup.scala 33:37]
  wire [3:0] _T_1574 = _T_433 ? 4'h2 : _T_1573; // @[Lookup.scala 33:37]
  wire [3:0] _T_1575 = _T_431 ? 4'h2 : _T_1574; // @[Lookup.scala 33:37]
  wire [3:0] _T_1576 = _T_429 ? 4'h2 : _T_1575; // @[Lookup.scala 33:37]
  wire [3:0] _T_1577 = _T_427 ? 4'h2 : _T_1576; // @[Lookup.scala 33:37]
  wire [3:0] _T_1578 = _T_425 ? 4'h2 : _T_1577; // @[Lookup.scala 33:37]
  wire [3:0] _T_1579 = _T_423 ? 4'h2 : _T_1578; // @[Lookup.scala 33:37]
  wire [3:0] _T_1580 = _T_421 ? 4'h2 : _T_1579; // @[Lookup.scala 33:37]
  wire [3:0] _T_1581 = _T_419 ? 4'h2 : _T_1580; // @[Lookup.scala 33:37]
  wire [3:0] _T_1582 = _T_417 ? 4'h2 : _T_1581; // @[Lookup.scala 33:37]
  wire [3:0] _T_1583 = _T_415 ? 4'h2 : _T_1582; // @[Lookup.scala 33:37]
  wire [3:0] _T_1584 = _T_413 ? 4'h2 : _T_1583; // @[Lookup.scala 33:37]
  wire [3:0] _T_1585 = _T_411 ? 4'h2 : _T_1584; // @[Lookup.scala 33:37]
  wire [3:0] _T_1586 = _T_409 ? 4'h2 : _T_1585; // @[Lookup.scala 33:37]
  wire [3:0] _T_1587 = _T_407 ? 4'h2 : _T_1586; // @[Lookup.scala 33:37]
  wire [3:0] _T_1588 = _T_405 ? 4'h2 : _T_1587; // @[Lookup.scala 33:37]
  wire [3:0] _T_1589 = _T_403 ? 4'h2 : _T_1588; // @[Lookup.scala 33:37]
  wire [3:0] _T_1590 = _T_401 ? 4'h2 : _T_1589; // @[Lookup.scala 33:37]
  wire [3:0] _T_1591 = _T_399 ? 4'h2 : _T_1590; // @[Lookup.scala 33:37]
  wire [3:0] _T_1592 = _T_397 ? 4'h2 : _T_1591; // @[Lookup.scala 33:37]
  wire [3:0] _T_1593 = _T_395 ? 4'h2 : _T_1592; // @[Lookup.scala 33:37]
  wire [3:0] _T_1594 = _T_393 ? 4'h2 : _T_1593; // @[Lookup.scala 33:37]
  wire [3:0] _T_1595 = _T_391 ? 4'h2 : _T_1594; // @[Lookup.scala 33:37]
  wire [3:0] _T_1596 = _T_389 ? 4'h2 : _T_1595; // @[Lookup.scala 33:37]
  wire [3:0] _T_1597 = _T_387 ? 4'h2 : _T_1596; // @[Lookup.scala 33:37]
  wire [3:0] _T_1598 = _T_385 ? 4'h2 : _T_1597; // @[Lookup.scala 33:37]
  wire [3:0] _T_1599 = _T_383 ? 4'h2 : _T_1598; // @[Lookup.scala 33:37]
  wire [3:0] _T_1600 = _T_381 ? 4'h2 : _T_1599; // @[Lookup.scala 33:37]
  wire [3:0] _T_1601 = _T_379 ? 4'h2 : _T_1600; // @[Lookup.scala 33:37]
  wire [3:0] _T_1602 = _T_377 ? 4'h2 : _T_1601; // @[Lookup.scala 33:37]
  wire [3:0] _T_1603 = _T_375 ? 4'h2 : _T_1602; // @[Lookup.scala 33:37]
  wire [3:0] _T_1604 = _T_373 ? 4'h2 : _T_1603; // @[Lookup.scala 33:37]
  wire [3:0] _T_1605 = _T_371 ? 4'h2 : _T_1604; // @[Lookup.scala 33:37]
  wire [3:0] _T_1606 = _T_369 ? 4'h2 : _T_1605; // @[Lookup.scala 33:37]
  wire [3:0] _T_1607 = _T_367 ? 4'h2 : _T_1606; // @[Lookup.scala 33:37]
  wire [3:0] _T_1608 = _T_365 ? 4'h2 : _T_1607; // @[Lookup.scala 33:37]
  wire [3:0] _T_1609 = _T_363 ? 4'h2 : _T_1608; // @[Lookup.scala 33:37]
  wire [3:0] _T_1610 = _T_361 ? 4'h2 : _T_1609; // @[Lookup.scala 33:37]
  wire [3:0] _T_1611 = _T_359 ? 4'h2 : _T_1610; // @[Lookup.scala 33:37]
  wire [3:0] _T_1612 = _T_357 ? 4'h2 : _T_1611; // @[Lookup.scala 33:37]
  wire [3:0] _T_1613 = _T_355 ? 4'h2 : _T_1612; // @[Lookup.scala 33:37]
  wire [3:0] _T_1614 = _T_353 ? 4'h2 : _T_1613; // @[Lookup.scala 33:37]
  wire [3:0] _T_1615 = _T_351 ? 4'h2 : _T_1614; // @[Lookup.scala 33:37]
  wire [3:0] _T_1616 = _T_349 ? 4'h2 : _T_1615; // @[Lookup.scala 33:37]
  wire [3:0] _T_1617 = _T_347 ? 4'h2 : _T_1616; // @[Lookup.scala 33:37]
  wire [3:0] _T_1618 = _T_345 ? 4'h2 : _T_1617; // @[Lookup.scala 33:37]
  wire [3:0] _T_1619 = _T_343 ? 4'h2 : _T_1618; // @[Lookup.scala 33:37]
  wire [3:0] _T_1620 = _T_341 ? 4'h2 : _T_1619; // @[Lookup.scala 33:37]
  wire [3:0] _T_1621 = _T_339 ? 4'h2 : _T_1620; // @[Lookup.scala 33:37]
  wire [3:0] _T_1622 = _T_337 ? 4'h2 : _T_1621; // @[Lookup.scala 33:37]
  wire [3:0] _T_1623 = _T_335 ? 4'h2 : _T_1622; // @[Lookup.scala 33:37]
  wire [3:0] _T_1624 = _T_333 ? 4'h2 : _T_1623; // @[Lookup.scala 33:37]
  wire [3:0] _T_1625 = _T_331 ? 4'h2 : _T_1624; // @[Lookup.scala 33:37]
  wire [3:0] _T_1626 = _T_329 ? 4'h2 : _T_1625; // @[Lookup.scala 33:37]
  wire [3:0] _T_1627 = _T_327 ? 4'h2 : _T_1626; // @[Lookup.scala 33:37]
  wire [3:0] _T_1628 = _T_325 ? 4'h2 : _T_1627; // @[Lookup.scala 33:37]
  wire [3:0] _T_1629 = _T_323 ? 4'h2 : _T_1628; // @[Lookup.scala 33:37]
  wire [3:0] _T_1630 = _T_321 ? 4'h2 : _T_1629; // @[Lookup.scala 33:37]
  wire [3:0] _T_1631 = _T_319 ? 4'h2 : _T_1630; // @[Lookup.scala 33:37]
  wire [3:0] _T_1632 = _T_317 ? 4'h2 : _T_1631; // @[Lookup.scala 33:37]
  wire [3:0] _T_1633 = _T_315 ? 4'h2 : _T_1632; // @[Lookup.scala 33:37]
  wire [3:0] _T_1634 = _T_313 ? 4'h2 : _T_1633; // @[Lookup.scala 33:37]
  wire [3:0] _T_1635 = _T_311 ? 4'h2 : _T_1634; // @[Lookup.scala 33:37]
  wire [3:0] _T_1636 = _T_309 ? 4'h2 : _T_1635; // @[Lookup.scala 33:37]
  wire [3:0] _T_1637 = _T_307 ? 4'h2 : _T_1636; // @[Lookup.scala 33:37]
  wire [3:0] _T_1638 = _T_305 ? 4'h2 : _T_1637; // @[Lookup.scala 33:37]
  wire [3:0] _T_1639 = _T_303 ? 4'h2 : _T_1638; // @[Lookup.scala 33:37]
  wire [3:0] _T_1640 = _T_301 ? 4'h2 : _T_1639; // @[Lookup.scala 33:37]
  wire [3:0] _T_1641 = _T_299 ? 4'h2 : _T_1640; // @[Lookup.scala 33:37]
  wire [3:0] _T_1642 = _T_297 ? 4'h2 : _T_1641; // @[Lookup.scala 33:37]
  wire [3:0] _T_1643 = _T_295 ? 4'h2 : _T_1642; // @[Lookup.scala 33:37]
  wire [3:0] _T_1644 = _T_293 ? 4'h2 : _T_1643; // @[Lookup.scala 33:37]
  wire [3:0] _T_1645 = _T_291 ? 4'h2 : _T_1644; // @[Lookup.scala 33:37]
  wire [3:0] _T_1646 = _T_289 ? 4'h2 : _T_1645; // @[Lookup.scala 33:37]
  wire [3:0] _T_1647 = _T_287 ? 4'h2 : _T_1646; // @[Lookup.scala 33:37]
  wire [3:0] _T_1648 = _T_285 ? 4'h2 : _T_1647; // @[Lookup.scala 33:37]
  wire [3:0] _T_1649 = _T_283 ? 4'h2 : _T_1648; // @[Lookup.scala 33:37]
  wire [3:0] _T_1650 = _T_281 ? 4'h2 : _T_1649; // @[Lookup.scala 33:37]
  wire [3:0] _T_1651 = _T_279 ? 4'h2 : _T_1650; // @[Lookup.scala 33:37]
  wire [3:0] _T_1652 = _T_277 ? 4'h2 : _T_1651; // @[Lookup.scala 33:37]
  wire [3:0] _T_1653 = _T_275 ? 4'h2 : _T_1652; // @[Lookup.scala 33:37]
  wire [3:0] _T_1654 = _T_273 ? 4'h2 : _T_1653; // @[Lookup.scala 33:37]
  wire [3:0] _T_1655 = _T_271 ? 4'h2 : _T_1654; // @[Lookup.scala 33:37]
  wire [3:0] _T_1656 = _T_269 ? 4'h2 : _T_1655; // @[Lookup.scala 33:37]
  wire [3:0] _T_1657 = _T_267 ? 4'h2 : _T_1656; // @[Lookup.scala 33:37]
  wire [3:0] _T_1658 = _T_265 ? 4'h2 : _T_1657; // @[Lookup.scala 33:37]
  wire [3:0] _T_1659 = _T_263 ? 4'h2 : _T_1658; // @[Lookup.scala 33:37]
  wire [3:0] _T_1660 = _T_261 ? 4'h2 : _T_1659; // @[Lookup.scala 33:37]
  wire [3:0] _T_1661 = _T_259 ? 4'h2 : _T_1660; // @[Lookup.scala 33:37]
  wire [3:0] _T_1662 = _T_257 ? 4'h2 : _T_1661; // @[Lookup.scala 33:37]
  wire [3:0] _T_1663 = _T_255 ? 4'h2 : _T_1662; // @[Lookup.scala 33:37]
  wire [3:0] _T_1664 = _T_253 ? 4'h2 : _T_1663; // @[Lookup.scala 33:37]
  wire [3:0] _T_1665 = _T_251 ? 4'h2 : _T_1664; // @[Lookup.scala 33:37]
  wire [3:0] _T_1666 = _T_249 ? 4'h2 : _T_1665; // @[Lookup.scala 33:37]
  wire [3:0] _T_1667 = _T_247 ? 4'h8 : _T_1666; // @[Lookup.scala 33:37]
  wire [3:0] _T_1668 = _T_245 ? 4'h1 : _T_1667; // @[Lookup.scala 33:37]
  wire [3:0] _T_1669 = _T_243 ? 4'h1 : _T_1668; // @[Lookup.scala 33:37]
  wire [3:0] _T_1670 = _T_241 ? 4'h1 : _T_1669; // @[Lookup.scala 33:37]
  wire [3:0] _T_1671 = _T_239 ? 4'h1 : _T_1670; // @[Lookup.scala 33:37]
  wire [3:0] _T_1672 = _T_237 ? 4'h1 : _T_1671; // @[Lookup.scala 33:37]
  wire [3:0] _T_1673 = _T_235 ? 4'h1 : _T_1672; // @[Lookup.scala 33:37]
  wire [3:0] _T_1674 = _T_233 ? 4'h4 : _T_1673; // @[Lookup.scala 33:37]
  wire [3:0] _T_1675 = _T_231 ? 4'h4 : _T_1674; // @[Lookup.scala 33:37]
  wire [3:0] _T_1676 = _T_229 ? 4'h4 : _T_1675; // @[Lookup.scala 33:37]
  wire [3:0] _T_1677 = _T_227 ? 4'h4 : _T_1676; // @[Lookup.scala 33:37]
  wire [3:0] _T_1678 = _T_225 ? 4'h4 : _T_1677; // @[Lookup.scala 33:37]
  wire [3:0] _T_1679 = _T_223 ? 4'h4 : _T_1678; // @[Lookup.scala 33:37]
  wire [3:0] _T_1680 = _T_221 ? 4'h4 : _T_1679; // @[Lookup.scala 33:37]
  wire [3:0] _T_1681 = _T_219 ? 4'h4 : _T_1680; // @[Lookup.scala 33:37]
  wire [3:0] _T_1682 = _T_217 ? 4'h4 : _T_1681; // @[Lookup.scala 33:37]
  wire [3:0] _T_1683 = _T_215 ? 4'h4 : _T_1682; // @[Lookup.scala 33:37]
  wire [3:0] _T_1684 = _T_213 ? 4'h4 : _T_1683; // @[Lookup.scala 33:37]
  wire [3:0] _T_1685 = _T_211 ? 4'h4 : _T_1684; // @[Lookup.scala 33:37]
  wire [3:0] _T_1686 = _T_209 ? 4'h4 : _T_1685; // @[Lookup.scala 33:37]
  wire [3:0] _T_1687 = _T_207 ? 4'h8 : _T_1686; // @[Lookup.scala 33:37]
  wire [3:0] _T_1688 = _T_205 ? 4'h1 : _T_1687; // @[Lookup.scala 33:37]
  wire [3:0] _T_1689 = _T_203 ? 4'h6 : _T_1688; // @[Lookup.scala 33:37]
  wire [3:0] _T_1690 = _T_201 ? 4'h8 : _T_1689; // @[Lookup.scala 33:37]
  wire [3:0] _T_1691 = _T_199 ? 4'h1 : _T_1690; // @[Lookup.scala 33:37]
  wire [3:0] _T_1692 = _T_197 ? 4'h1 : _T_1691; // @[Lookup.scala 33:37]
  wire [3:0] _T_1693 = _T_195 ? 4'h1 : _T_1692; // @[Lookup.scala 33:37]
  wire [3:0] _T_1694 = _T_193 ? 4'h4 : _T_1693; // @[Lookup.scala 33:37]
  wire [3:0] _T_1695 = _T_191 ? 4'h4 : _T_1694; // @[Lookup.scala 33:37]
  wire [3:0] _T_1696 = _T_189 ? 4'h6 : _T_1695; // @[Lookup.scala 33:37]
  wire [3:0] _T_1697 = _T_187 ? 4'h0 : _T_1696; // @[Lookup.scala 33:37]
  wire [3:0] _T_1698 = _T_185 ? 4'h1 : _T_1697; // @[Lookup.scala 33:37]
  wire [3:0] _T_1699 = _T_183 ? 4'h6 : _T_1698; // @[Lookup.scala 33:37]
  wire [3:0] _T_1700 = _T_181 ? 4'h0 : _T_1699; // @[Lookup.scala 33:37]
  wire [3:0] _T_1701 = _T_179 ? 4'h4 : _T_1700; // @[Lookup.scala 33:37]
  wire [3:0] _T_1702 = _T_177 ? 4'h4 : _T_1701; // @[Lookup.scala 33:37]
  wire [3:0] _T_1703 = _T_175 ? 4'h6 : _T_1702; // @[Lookup.scala 33:37]
  wire [3:0] _T_1704 = _T_173 ? 4'h0 : _T_1703; // @[Lookup.scala 33:37]
  wire [3:0] _T_1705 = _T_171 ? 4'h0 : _T_1704; // @[Lookup.scala 33:37]
  wire [3:0] _T_1706 = _T_169 ? 4'h0 : _T_1705; // @[Lookup.scala 33:37]
  wire [3:0] _T_1707 = _T_167 ? 4'h6 : _T_1706; // @[Lookup.scala 33:37]
  wire [3:0] _T_1708 = _T_165 ? 4'h6 : _T_1707; // @[Lookup.scala 33:37]
  wire [3:0] _T_1709 = _T_163 ? 4'h6 : _T_1708; // @[Lookup.scala 33:37]
  wire [3:0] _T_1710 = _T_161 ? 4'h6 : _T_1709; // @[Lookup.scala 33:37]
  wire [3:0] _T_1711 = _T_159 ? 4'h6 : _T_1710; // @[Lookup.scala 33:37]
  wire [3:0] _T_1712 = _T_157 ? 4'h6 : _T_1711; // @[Lookup.scala 33:37]
  wire [3:0] _T_1713 = _T_155 ? 4'h6 : _T_1712; // @[Lookup.scala 33:37]
  wire [3:0] _T_1714 = _T_153 ? 4'h6 : _T_1713; // @[Lookup.scala 33:37]
  wire [3:0] _T_1715 = _T_151 ? 4'h6 : _T_1714; // @[Lookup.scala 33:37]
  wire [3:0] _T_1716 = _T_149 ? 4'h6 : _T_1715; // @[Lookup.scala 33:37]
  wire [3:0] _T_1717 = _T_147 ? 4'h6 : _T_1716; // @[Lookup.scala 33:37]
  wire [3:0] _T_1718 = _T_145 ? 4'h6 : _T_1717; // @[Lookup.scala 33:37]
  wire [3:0] _T_1719 = _T_143 ? 4'h6 : _T_1718; // @[Lookup.scala 33:37]
  wire [3:0] _T_1720 = _T_141 ? 4'h6 : _T_1719; // @[Lookup.scala 33:37]
  wire [3:0] _T_1721 = _T_139 ? 4'h6 : _T_1720; // @[Lookup.scala 33:37]
  wire [3:0] _T_1722 = _T_137 ? 4'h4 : _T_1721; // @[Lookup.scala 33:37]
  wire [3:0] _T_1723 = _T_135 ? 4'h4 : _T_1722; // @[Lookup.scala 33:37]
  wire [3:0] _T_1724 = _T_133 ? 4'h4 : _T_1723; // @[Lookup.scala 33:37]
  wire [3:0] _T_1725 = _T_131 ? 4'h4 : _T_1724; // @[Lookup.scala 33:37]
  wire [3:0] _T_1726 = _T_129 ? 4'h6 : _T_1725; // @[Lookup.scala 33:37]
  wire [3:0] _T_1727 = _T_127 ? 4'h1 : _T_1726; // @[Lookup.scala 33:37]
  wire [3:0] _T_1728 = _T_125 ? 4'h5 : _T_1727; // @[Lookup.scala 33:37]
  wire [3:0] _T_1729 = _T_123 ? 4'h5 : _T_1728; // @[Lookup.scala 33:37]
  wire [3:0] _T_1730 = _T_121 ? 4'h5 : _T_1729; // @[Lookup.scala 33:37]
  wire [3:0] _T_1731 = _T_119 ? 4'h5 : _T_1730; // @[Lookup.scala 33:37]
  wire [3:0] _T_1732 = _T_117 ? 4'h5 : _T_1731; // @[Lookup.scala 33:37]
  wire [3:0] _T_1733 = _T_115 ? 4'h5 : _T_1732; // @[Lookup.scala 33:37]
  wire [3:0] _T_1734 = _T_113 ? 4'h5 : _T_1733; // @[Lookup.scala 33:37]
  wire [3:0] _T_1735 = _T_111 ? 4'h5 : _T_1734; // @[Lookup.scala 33:37]
  wire [3:0] _T_1736 = _T_109 ? 4'h5 : _T_1735; // @[Lookup.scala 33:37]
  wire [3:0] _T_1737 = _T_107 ? 4'h5 : _T_1736; // @[Lookup.scala 33:37]
  wire [3:0] _T_1738 = _T_105 ? 4'h5 : _T_1737; // @[Lookup.scala 33:37]
  wire [3:0] _T_1739 = _T_103 ? 4'h5 : _T_1738; // @[Lookup.scala 33:37]
  wire [3:0] _T_1740 = _T_101 ? 4'h5 : _T_1739; // @[Lookup.scala 33:37]
  wire [3:0] _T_1741 = _T_99 ? 4'h1 : _T_1740; // @[Lookup.scala 33:37]
  wire [3:0] _T_1742 = _T_97 ? 4'h4 : _T_1741; // @[Lookup.scala 33:37]
  wire [3:0] _T_1743 = _T_95 ? 4'h4 : _T_1742; // @[Lookup.scala 33:37]
  wire [3:0] _T_1744 = _T_93 ? 4'h4 : _T_1743; // @[Lookup.scala 33:37]
  wire [3:0] _T_1745 = _T_91 ? 4'h6 : _T_1744; // @[Lookup.scala 33:37]
  wire [3:0] _T_1746 = _T_89 ? 4'h6 : _T_1745; // @[Lookup.scala 33:37]
  wire [3:0] _T_1747 = _T_87 ? 4'h6 : _T_1746; // @[Lookup.scala 33:37]
  wire [3:0] _T_1748 = _T_85 ? 4'h6 : _T_1747; // @[Lookup.scala 33:37]
  wire [3:0] _T_1749 = _T_83 ? 4'h6 : _T_1748; // @[Lookup.scala 33:37]
  wire [3:0] _T_1750 = _T_81 ? 4'h6 : _T_1749; // @[Lookup.scala 33:37]
  wire [3:0] _T_1751 = _T_79 ? 4'h6 : _T_1750; // @[Lookup.scala 33:37]
  wire [3:0] _T_1752 = _T_77 ? 4'h6 : _T_1751; // @[Lookup.scala 33:37]
  wire [3:0] _T_1753 = _T_75 ? 4'h6 : _T_1752; // @[Lookup.scala 33:37]
  wire [3:0] _T_1754 = _T_73 ? 4'h4 : _T_1753; // @[Lookup.scala 33:37]
  wire [3:0] _T_1755 = _T_71 ? 4'h4 : _T_1754; // @[Lookup.scala 33:37]
  wire [3:0] _T_1756 = _T_69 ? 4'h4 : _T_1755; // @[Lookup.scala 33:37]
  wire [3:0] _T_1757 = _T_67 ? 4'h4 : _T_1756; // @[Lookup.scala 33:37]
  wire [3:0] _T_1758 = _T_65 ? 4'h4 : _T_1757; // @[Lookup.scala 33:37]
  wire [3:0] _T_1759 = _T_63 ? 4'h4 : _T_1758; // @[Lookup.scala 33:37]
  wire [3:0] _T_1760 = _T_61 ? 4'h4 : _T_1759; // @[Lookup.scala 33:37]
  wire [3:0] _T_1761 = _T_59 ? 4'h4 : _T_1760; // @[Lookup.scala 33:37]
  wire [3:0] _T_1762 = _T_57 ? 4'h0 : _T_1761; // @[Lookup.scala 33:37]
  wire [3:0] _T_1763 = _T_55 ? 4'h0 : _T_1762; // @[Lookup.scala 33:37]
  wire [3:0] _T_1764 = _T_53 ? 4'h0 : _T_1763; // @[Lookup.scala 33:37]
  wire [3:0] _T_1765 = _T_51 ? 4'h0 : _T_1764; // @[Lookup.scala 33:37]
  wire [3:0] _T_1766 = _T_49 ? 4'h0 : _T_1765; // @[Lookup.scala 33:37]
  wire [3:0] _T_1767 = _T_47 ? 4'h0 : _T_1766; // @[Lookup.scala 33:37]
  wire [3:0] _T_1768 = _T_45 ? 4'h0 : _T_1767; // @[Lookup.scala 33:37]
  wire [3:0] _T_1769 = _T_43 ? 4'h0 : _T_1768; // @[Lookup.scala 33:37]
  wire [3:0] _T_1770 = _T_41 ? 4'h6 : _T_1769; // @[Lookup.scala 33:37]
  wire [3:0] _T_1771 = _T_39 ? 4'h6 : _T_1770; // @[Lookup.scala 33:37]
  wire [3:0] _T_1772 = _T_37 ? 4'h6 : _T_1771; // @[Lookup.scala 33:37]
  wire [3:0] _T_1773 = _T_35 ? 4'h6 : _T_1772; // @[Lookup.scala 33:37]
  wire [3:0] _T_1774 = _T_33 ? 4'h6 : _T_1773; // @[Lookup.scala 33:37]
  wire [3:0] _T_1775 = _T_31 ? 4'h6 : _T_1774; // @[Lookup.scala 33:37]
  wire [3:0] _T_1776 = _T_29 ? 4'h6 : _T_1775; // @[Lookup.scala 33:37]
  wire [3:0] _T_1777 = _T_27 ? 4'h6 : _T_1776; // @[Lookup.scala 33:37]
  wire [3:0] _T_1778 = _T_25 ? 4'h6 : _T_1777; // @[Lookup.scala 33:37]
  wire [3:0] _T_1779 = _T_23 ? 4'h6 : _T_1778; // @[Lookup.scala 33:37]
  wire [3:0] _T_1780 = _T_21 ? 4'h6 : _T_1779; // @[Lookup.scala 33:37]
  wire [3:0] _T_1781 = _T_19 ? 4'h6 : _T_1780; // @[Lookup.scala 33:37]
  wire [3:0] _T_1782 = _T_17 ? 4'h6 : _T_1781; // @[Lookup.scala 33:37]
  wire [3:0] _T_1783 = _T_15 ? 4'h6 : _T_1782; // @[Lookup.scala 33:37]
  wire [3:0] _T_1784 = _T_13 ? 4'h6 : _T_1783; // @[Lookup.scala 33:37]
  wire [3:0] _T_1785 = _T_11 ? 4'h6 : _T_1784; // @[Lookup.scala 33:37]
  wire [3:0] _T_1786 = _T_9 ? 4'h6 : _T_1785; // @[Lookup.scala 33:37]
  wire [3:0] _T_1787 = _T_7 ? 4'h6 : _T_1786; // @[Lookup.scala 33:37]
  wire [3:0] _T_1788 = _T_5 ? 4'h6 : _T_1787; // @[Lookup.scala 33:37]
  wire [3:0] _T_1789 = _T_3 ? 4'h6 : _T_1788; // @[Lookup.scala 33:37]
  wire [3:0] decodeList_1 = _T_1 ? 4'h6 : _T_1789; // @[Lookup.scala 33:37]
  wire [5:0] _T_1790 = _T_895 ? 6'h3e : 6'h0; // @[Lookup.scala 33:37]
  wire [5:0] _T_1791 = _T_893 ? 6'h36 : _T_1790; // @[Lookup.scala 33:37]
  wire [5:0] _T_1792 = _T_891 ? 6'h2e : _T_1791; // @[Lookup.scala 33:37]
  wire [5:0] _T_1793 = _T_889 ? 6'h27 : _T_1792; // @[Lookup.scala 33:37]
  wire [5:0] _T_1794 = _T_887 ? 6'h26 : _T_1793; // @[Lookup.scala 33:37]
  wire [5:0] _T_1795 = _T_885 ? 6'h25 : _T_1794; // @[Lookup.scala 33:37]
  wire [5:0] _T_1796 = _T_883 ? 6'h3d : _T_1795; // @[Lookup.scala 33:37]
  wire [5:0] _T_1797 = _T_881 ? 6'h35 : _T_1796; // @[Lookup.scala 33:37]
  wire [5:0] _T_1798 = _T_879 ? 6'h2d : _T_1797; // @[Lookup.scala 33:37]
  wire [6:0] _T_1799 = _T_877 ? 7'h7c : {{1'd0}, _T_1798}; // @[Lookup.scala 33:37]
  wire [6:0] _T_1800 = _T_875 ? 7'h74 : _T_1799; // @[Lookup.scala 33:37]
  wire [6:0] _T_1801 = _T_873 ? 7'h6c : _T_1800; // @[Lookup.scala 33:37]
  wire [6:0] _T_1802 = _T_871 ? 7'h63 : _T_1801; // @[Lookup.scala 33:37]
  wire [6:0] _T_1803 = _T_869 ? 7'h62 : _T_1802; // @[Lookup.scala 33:37]
  wire [6:0] _T_1804 = _T_867 ? 7'h79 : _T_1803; // @[Lookup.scala 33:37]
  wire [6:0] _T_1805 = _T_865 ? 7'h71 : _T_1804; // @[Lookup.scala 33:37]
  wire [6:0] _T_1806 = _T_863 ? 7'h69 : _T_1805; // @[Lookup.scala 33:37]
  wire [6:0] _T_1807 = _T_861 ? 7'h5e : _T_1806; // @[Lookup.scala 33:37]
  wire [6:0] _T_1808 = _T_859 ? 7'h56 : _T_1807; // @[Lookup.scala 33:37]
  wire [6:0] _T_1809 = _T_857 ? 7'h4e : _T_1808; // @[Lookup.scala 33:37]
  wire [6:0] _T_1810 = _T_855 ? 7'h46 : _T_1809; // @[Lookup.scala 33:37]
  wire [6:0] _T_1811 = _T_853 ? 7'h55 : _T_1810; // @[Lookup.scala 33:37]
  wire [6:0] _T_1812 = _T_851 ? 7'h4d : _T_1811; // @[Lookup.scala 33:37]
  wire [6:0] _T_1813 = _T_849 ? 7'h45 : _T_1812; // @[Lookup.scala 33:37]
  wire [6:0] _T_1814 = _T_847 ? 7'h54 : _T_1813; // @[Lookup.scala 33:37]
  wire [6:0] _T_1815 = _T_845 ? 7'h4c : _T_1814; // @[Lookup.scala 33:37]
  wire [6:0] _T_1816 = _T_843 ? 7'h44 : _T_1815; // @[Lookup.scala 33:37]
  wire [6:0] _T_1817 = _T_841 ? 7'h5b : _T_1816; // @[Lookup.scala 33:37]
  wire [6:0] _T_1818 = _T_839 ? 7'h53 : _T_1817; // @[Lookup.scala 33:37]
  wire [6:0] _T_1819 = _T_837 ? 7'h4b : _T_1818; // @[Lookup.scala 33:37]
  wire [6:0] _T_1820 = _T_835 ? 7'h43 : _T_1819; // @[Lookup.scala 33:37]
  wire [6:0] _T_1821 = _T_833 ? 7'h5a : _T_1820; // @[Lookup.scala 33:37]
  wire [6:0] _T_1822 = _T_831 ? 7'h52 : _T_1821; // @[Lookup.scala 33:37]
  wire [6:0] _T_1823 = _T_829 ? 7'h4a : _T_1822; // @[Lookup.scala 33:37]
  wire [6:0] _T_1824 = _T_827 ? 7'h42 : _T_1823; // @[Lookup.scala 33:37]
  wire [6:0] _T_1825 = _T_825 ? 7'h66 : _T_1824; // @[Lookup.scala 33:37]
  wire [6:0] _T_1826 = _T_823 ? 7'h65 : _T_1825; // @[Lookup.scala 33:37]
  wire [6:0] _T_1827 = _T_821 ? 7'h64 : _T_1826; // @[Lookup.scala 33:37]
  wire [6:0] _T_1828 = _T_819 ? 7'h27 : _T_1827; // @[Lookup.scala 33:37]
  wire [6:0] _T_1829 = _T_817 ? 7'h26 : _T_1828; // @[Lookup.scala 33:37]
  wire [6:0] _T_1830 = _T_815 ? 7'h3e : _T_1829; // @[Lookup.scala 33:37]
  wire [6:0] _T_1831 = _T_813 ? 7'h36 : _T_1830; // @[Lookup.scala 33:37]
  wire [6:0] _T_1832 = _T_811 ? 7'h2e : _T_1831; // @[Lookup.scala 33:37]
  wire [6:0] _T_1833 = _T_809 ? 7'h25 : _T_1832; // @[Lookup.scala 33:37]
  wire [6:0] _T_1834 = _T_807 ? 7'h24 : _T_1833; // @[Lookup.scala 33:37]
  wire [6:0] _T_1835 = _T_805 ? 7'h3d : _T_1834; // @[Lookup.scala 33:37]
  wire [6:0] _T_1836 = _T_803 ? 7'h35 : _T_1835; // @[Lookup.scala 33:37]
  wire [6:0] _T_1837 = _T_801 ? 7'h2d : _T_1836; // @[Lookup.scala 33:37]
  wire [6:0] _T_1838 = _T_799 ? 7'h7f : _T_1837; // @[Lookup.scala 33:37]
  wire [6:0] _T_1839 = _T_797 ? 7'h77 : _T_1838; // @[Lookup.scala 33:37]
  wire [6:0] _T_1840 = _T_795 ? 7'h6f : _T_1839; // @[Lookup.scala 33:37]
  wire [6:0] _T_1841 = _T_793 ? 7'h67 : _T_1840; // @[Lookup.scala 33:37]
  wire [6:0] _T_1842 = _T_791 ? 7'h3b : _T_1841; // @[Lookup.scala 33:37]
  wire [6:0] _T_1843 = _T_789 ? 7'h33 : _T_1842; // @[Lookup.scala 33:37]
  wire [6:0] _T_1844 = _T_787 ? 7'h2b : _T_1843; // @[Lookup.scala 33:37]
  wire [6:0] _T_1845 = _T_785 ? 7'h23 : _T_1844; // @[Lookup.scala 33:37]
  wire [6:0] _T_1846 = _T_783 ? 7'h29 : _T_1845; // @[Lookup.scala 33:37]
  wire [6:0] _T_1847 = _T_781 ? 7'h21 : _T_1846; // @[Lookup.scala 33:37]
  wire [6:0] _T_1848 = _T_779 ? 7'h38 : _T_1847; // @[Lookup.scala 33:37]
  wire [6:0] _T_1849 = _T_777 ? 7'h30 : _T_1848; // @[Lookup.scala 33:37]
  wire [6:0] _T_1850 = _T_775 ? 7'h35 : _T_1849; // @[Lookup.scala 33:37]
  wire [6:0] _T_1851 = _T_773 ? 7'h3b : _T_1850; // @[Lookup.scala 33:37]
  wire [6:0] _T_1852 = _T_771 ? 7'h24 : _T_1851; // @[Lookup.scala 33:37]
  wire [6:0] _T_1853 = _T_769 ? 7'h4 : _T_1852; // @[Lookup.scala 33:37]
  wire [6:0] _T_1854 = _T_767 ? 7'h5 : _T_1853; // @[Lookup.scala 33:37]
  wire [6:0] _T_1855 = _T_765 ? 7'h5 : _T_1854; // @[Lookup.scala 33:37]
  wire [6:0] _T_1856 = _T_763 ? 7'h56 : _T_1855; // @[Lookup.scala 33:37]
  wire [6:0] _T_1857 = _T_761 ? 7'h3c : _T_1856; // @[Lookup.scala 33:37]
  wire [6:0] _T_1858 = _T_759 ? 7'h34 : _T_1857; // @[Lookup.scala 33:37]
  wire [6:0] _T_1859 = _T_757 ? 7'h2c : _T_1858; // @[Lookup.scala 33:37]
  wire [6:0] _T_1860 = _T_755 ? 7'h1d : _T_1859; // @[Lookup.scala 33:37]
  wire [6:0] _T_1861 = _T_753 ? 7'h1c : _T_1860; // @[Lookup.scala 33:37]
  wire [6:0] _T_1862 = _T_751 ? 7'h14 : _T_1861; // @[Lookup.scala 33:37]
  wire [6:0] _T_1863 = _T_749 ? 7'hc : _T_1862; // @[Lookup.scala 33:37]
  wire [6:0] _T_1864 = _T_747 ? 7'h7d : _T_1863; // @[Lookup.scala 33:37]
  wire [6:0] _T_1865 = _T_745 ? 7'h75 : _T_1864; // @[Lookup.scala 33:37]
  wire [6:0] _T_1866 = _T_743 ? 7'h6d : _T_1865; // @[Lookup.scala 33:37]
  wire [6:0] _T_1867 = _T_741 ? 7'h7e : _T_1866; // @[Lookup.scala 33:37]
  wire [6:0] _T_1868 = _T_739 ? 7'h76 : _T_1867; // @[Lookup.scala 33:37]
  wire [6:0] _T_1869 = _T_737 ? 7'h6e : _T_1868; // @[Lookup.scala 33:37]
  wire [6:0] _T_1870 = _T_735 ? 7'h70 : _T_1869; // @[Lookup.scala 33:37]
  wire [6:0] _T_1871 = _T_733 ? 7'h78 : _T_1870; // @[Lookup.scala 33:37]
  wire [6:0] _T_1872 = _T_731 ? 7'h15 : _T_1871; // @[Lookup.scala 33:37]
  wire [6:0] _T_1873 = _T_729 ? 7'hd : _T_1872; // @[Lookup.scala 33:37]
  wire [6:0] _T_1874 = _T_727 ? 7'h5 : _T_1873; // @[Lookup.scala 33:37]
  wire [6:0] _T_1875 = _T_725 ? 7'h16 : _T_1874; // @[Lookup.scala 33:37]
  wire [6:0] _T_1876 = _T_723 ? 7'he : _T_1875; // @[Lookup.scala 33:37]
  wire [6:0] _T_1877 = _T_721 ? 7'h6 : _T_1876; // @[Lookup.scala 33:37]
  wire [6:0] _T_1878 = _T_719 ? 7'h2f : _T_1877; // @[Lookup.scala 33:37]
  wire [6:0] _T_1879 = _T_717 ? 7'h3c : _T_1878; // @[Lookup.scala 33:37]
  wire [6:0] _T_1880 = _T_715 ? 7'h34 : _T_1879; // @[Lookup.scala 33:37]
  wire [6:0] _T_1881 = _T_713 ? 7'h2c : _T_1880; // @[Lookup.scala 33:37]
  wire [6:0] _T_1882 = _T_711 ? 7'h1d : _T_1881; // @[Lookup.scala 33:37]
  wire [6:0] _T_1883 = _T_709 ? 7'h1c : _T_1882; // @[Lookup.scala 33:37]
  wire [6:0] _T_1884 = _T_707 ? 7'h14 : _T_1883; // @[Lookup.scala 33:37]
  wire [6:0] _T_1885 = _T_705 ? 7'hc : _T_1884; // @[Lookup.scala 33:37]
  wire [6:0] _T_1886 = _T_703 ? 7'h4 : _T_1885; // @[Lookup.scala 33:37]
  wire [6:0] _T_1887 = _T_701 ? 7'h5f : _T_1886; // @[Lookup.scala 33:37]
  wire [6:0] _T_1888 = _T_699 ? 7'h57 : _T_1887; // @[Lookup.scala 33:37]
  wire [6:0] _T_1889 = _T_697 ? 7'h4f : _T_1888; // @[Lookup.scala 33:37]
  wire [6:0] _T_1890 = _T_695 ? 7'h47 : _T_1889; // @[Lookup.scala 33:37]
  wire [6:0] _T_1891 = _T_693 ? 7'h3a : _T_1890; // @[Lookup.scala 33:37]
  wire [6:0] _T_1892 = _T_691 ? 7'h32 : _T_1891; // @[Lookup.scala 33:37]
  wire [6:0] _T_1893 = _T_689 ? 7'h2a : _T_1892; // @[Lookup.scala 33:37]
  wire [6:0] _T_1894 = _T_687 ? 7'h22 : _T_1893; // @[Lookup.scala 33:37]
  wire [6:0] _T_1895 = _T_685 ? 7'h39 : _T_1894; // @[Lookup.scala 33:37]
  wire [6:0] _T_1896 = _T_683 ? 7'h31 : _T_1895; // @[Lookup.scala 33:37]
  wire [6:0] _T_1897 = _T_681 ? 7'h28 : _T_1896; // @[Lookup.scala 33:37]
  wire [6:0] _T_1898 = _T_679 ? 7'h20 : _T_1897; // @[Lookup.scala 33:37]
  wire [6:0] _T_1899 = _T_677 ? 7'h4f : _T_1898; // @[Lookup.scala 33:37]
  wire [6:0] _T_1900 = _T_675 ? 7'h47 : _T_1899; // @[Lookup.scala 33:37]
  wire [6:0] _T_1901 = _T_673 ? 7'h5d : _T_1900; // @[Lookup.scala 33:37]
  wire [6:0] _T_1902 = _T_671 ? 7'h55 : _T_1901; // @[Lookup.scala 33:37]
  wire [6:0] _T_1903 = _T_669 ? 7'h5c : _T_1902; // @[Lookup.scala 33:37]
  wire [6:0] _T_1904 = _T_667 ? 7'h54 : _T_1903; // @[Lookup.scala 33:37]
  wire [6:0] _T_1905 = _T_665 ? 7'h4b : _T_1904; // @[Lookup.scala 33:37]
  wire [6:0] _T_1906 = _T_663 ? 7'h43 : _T_1905; // @[Lookup.scala 33:37]
  wire [6:0] _T_1907 = _T_661 ? 7'h59 : _T_1906; // @[Lookup.scala 33:37]
  wire [6:0] _T_1908 = _T_659 ? 7'h51 : _T_1907; // @[Lookup.scala 33:37]
  wire [6:0] _T_1909 = _T_657 ? 7'h58 : _T_1908; // @[Lookup.scala 33:37]
  wire [6:0] _T_1910 = _T_655 ? 7'h50 : _T_1909; // @[Lookup.scala 33:37]
  wire [6:0] _T_1911 = _T_653 ? 7'h1a : _T_1910; // @[Lookup.scala 33:37]
  wire [6:0] _T_1912 = _T_651 ? 7'h56 : _T_1911; // @[Lookup.scala 33:37]
  wire [6:0] _T_1913 = _T_649 ? 7'h6f : _T_1912; // @[Lookup.scala 33:37]
  wire [6:0] _T_1914 = _T_647 ? 7'h74 : _T_1913; // @[Lookup.scala 33:37]
  wire [6:0] _T_1915 = _T_645 ? 7'h6a : _T_1914; // @[Lookup.scala 33:37]
  wire [6:0] _T_1916 = _T_643 ? 7'h1b : _T_1915; // @[Lookup.scala 33:37]
  wire [6:0] _T_1917 = _T_641 ? 7'h57 : _T_1916; // @[Lookup.scala 33:37]
  wire [6:0] _T_1918 = _T_639 ? 7'h57 : _T_1917; // @[Lookup.scala 33:37]
  wire [6:0] _T_1919 = _T_637 ? 7'h7a : _T_1918; // @[Lookup.scala 33:37]
  wire [6:0] _T_1920 = _T_635 ? 7'h72 : _T_1919; // @[Lookup.scala 33:37]
  wire [6:0] _T_1921 = _T_633 ? 7'h56 : _T_1920; // @[Lookup.scala 33:37]
  wire [6:0] _T_1922 = _T_631 ? 7'h56 : _T_1921; // @[Lookup.scala 33:37]
  wire [6:0] _T_1923 = _T_629 ? 7'h56 : _T_1922; // @[Lookup.scala 33:37]
  wire [6:0] _T_1924 = _T_627 ? 7'h56 : _T_1923; // @[Lookup.scala 33:37]
  wire [6:0] _T_1925 = _T_625 ? 7'h56 : _T_1924; // @[Lookup.scala 33:37]
  wire [6:0] _T_1926 = _T_623 ? 7'h56 : _T_1925; // @[Lookup.scala 33:37]
  wire [6:0] _T_1927 = _T_621 ? 7'h56 : _T_1926; // @[Lookup.scala 33:37]
  wire [6:0] _T_1928 = _T_619 ? 7'h56 : _T_1927; // @[Lookup.scala 33:37]
  wire [6:0] _T_1929 = _T_617 ? 7'h56 : _T_1928; // @[Lookup.scala 33:37]
  wire [6:0] _T_1930 = _T_615 ? 7'h56 : _T_1929; // @[Lookup.scala 33:37]
  wire [6:0] _T_1931 = _T_613 ? 7'h56 : _T_1930; // @[Lookup.scala 33:37]
  wire [6:0] _T_1932 = _T_611 ? 7'h57 : _T_1931; // @[Lookup.scala 33:37]
  wire [6:0] _T_1933 = _T_609 ? 7'h57 : _T_1932; // @[Lookup.scala 33:37]
  wire [6:0] _T_1934 = _T_607 ? 7'h57 : _T_1933; // @[Lookup.scala 33:37]
  wire [6:0] _T_1935 = _T_605 ? 7'h57 : _T_1934; // @[Lookup.scala 33:37]
  wire [6:0] _T_1936 = _T_603 ? 7'h56 : _T_1935; // @[Lookup.scala 33:37]
  wire [6:0] _T_1937 = _T_601 ? 7'h56 : _T_1936; // @[Lookup.scala 33:37]
  wire [6:0] _T_1938 = _T_599 ? 7'h56 : _T_1937; // @[Lookup.scala 33:37]
  wire [6:0] _T_1939 = _T_597 ? 7'h56 : _T_1938; // @[Lookup.scala 33:37]
  wire [6:0] _T_1940 = _T_595 ? 7'h46 : _T_1939; // @[Lookup.scala 33:37]
  wire [6:0] _T_1941 = _T_593 ? 7'h46 : _T_1940; // @[Lookup.scala 33:37]
  wire [6:0] _T_1942 = _T_591 ? 7'h42 : _T_1941; // @[Lookup.scala 33:37]
  wire [6:0] _T_1943 = _T_589 ? 7'h42 : _T_1942; // @[Lookup.scala 33:37]
  wire [6:0] _T_1944 = _T_587 ? 7'h42 : _T_1943; // @[Lookup.scala 33:37]
  wire [6:0] _T_1945 = _T_585 ? 7'h3a : _T_1944; // @[Lookup.scala 33:37]
  wire [6:0] _T_1946 = _T_583 ? 7'h41 : _T_1945; // @[Lookup.scala 33:37]
  wire [6:0] _T_1947 = _T_581 ? 7'h39 : _T_1946; // @[Lookup.scala 33:37]
  wire [6:0] _T_1948 = _T_579 ? 7'h40 : _T_1947; // @[Lookup.scala 33:37]
  wire [6:0] _T_1949 = _T_577 ? 7'h38 : _T_1948; // @[Lookup.scala 33:37]
  wire [6:0] _T_1950 = _T_575 ? 7'h3e : _T_1949; // @[Lookup.scala 33:37]
  wire [6:0] _T_1951 = _T_573 ? 7'h3e : _T_1950; // @[Lookup.scala 33:37]
  wire [6:0] _T_1952 = _T_571 ? 7'h3d : _T_1951; // @[Lookup.scala 33:37]
  wire [6:0] _T_1953 = _T_569 ? 7'h3d : _T_1952; // @[Lookup.scala 33:37]
  wire [6:0] _T_1954 = _T_567 ? 7'h3c : _T_1953; // @[Lookup.scala 33:37]
  wire [6:0] _T_1955 = _T_565 ? 7'h3c : _T_1954; // @[Lookup.scala 33:37]
  wire [6:0] _T_1956 = _T_563 ? 7'h3a : _T_1955; // @[Lookup.scala 33:37]
  wire [6:0] _T_1957 = _T_561 ? 7'h3a : _T_1956; // @[Lookup.scala 33:37]
  wire [6:0] _T_1958 = _T_559 ? 7'h39 : _T_1957; // @[Lookup.scala 33:37]
  wire [6:0] _T_1959 = _T_557 ? 7'h39 : _T_1958; // @[Lookup.scala 33:37]
  wire [6:0] _T_1960 = _T_555 ? 7'h38 : _T_1959; // @[Lookup.scala 33:37]
  wire [6:0] _T_1961 = _T_553 ? 7'h38 : _T_1960; // @[Lookup.scala 33:37]
  wire [6:0] _T_1962 = _T_551 ? 7'h1f : _T_1961; // @[Lookup.scala 33:37]
  wire [6:0] _T_1963 = _T_549 ? 7'hf : _T_1962; // @[Lookup.scala 33:37]
  wire [6:0] _T_1964 = _T_547 ? 7'h51 : _T_1963; // @[Lookup.scala 33:37]
  wire [6:0] _T_1965 = _T_545 ? 7'h50 : _T_1964; // @[Lookup.scala 33:37]
  wire [6:0] _T_1966 = _T_543 ? 7'h49 : _T_1965; // @[Lookup.scala 33:37]
  wire [6:0] _T_1967 = _T_541 ? 7'h48 : _T_1966; // @[Lookup.scala 33:37]
  wire [6:0] _T_1968 = _T_539 ? 7'h73 : _T_1967; // @[Lookup.scala 33:37]
  wire [6:0] _T_1969 = _T_537 ? 7'h6b : _T_1968; // @[Lookup.scala 33:37]
  wire [6:0] _T_1970 = _T_535 ? 7'h63 : _T_1969; // @[Lookup.scala 33:37]
  wire [6:0] _T_1971 = _T_533 ? 7'h5b : _T_1970; // @[Lookup.scala 33:37]
  wire [6:0] _T_1972 = _T_531 ? 7'h7b : _T_1971; // @[Lookup.scala 33:37]
  wire [6:0] _T_1973 = _T_529 ? 7'h72 : _T_1972; // @[Lookup.scala 33:37]
  wire [6:0] _T_1974 = _T_527 ? 7'h6a : _T_1973; // @[Lookup.scala 33:37]
  wire [6:0] _T_1975 = _T_525 ? 7'h62 : _T_1974; // @[Lookup.scala 33:37]
  wire [6:0] _T_1976 = _T_523 ? 7'h5a : _T_1975; // @[Lookup.scala 33:37]
  wire [6:0] _T_1977 = _T_521 ? 7'h7a : _T_1976; // @[Lookup.scala 33:37]
  wire [6:0] _T_1978 = _T_519 ? 7'h71 : _T_1977; // @[Lookup.scala 33:37]
  wire [6:0] _T_1979 = _T_517 ? 7'h69 : _T_1978; // @[Lookup.scala 33:37]
  wire [6:0] _T_1980 = _T_515 ? 7'h61 : _T_1979; // @[Lookup.scala 33:37]
  wire [6:0] _T_1981 = _T_513 ? 7'h59 : _T_1980; // @[Lookup.scala 33:37]
  wire [6:0] _T_1982 = _T_511 ? 7'h79 : _T_1981; // @[Lookup.scala 33:37]
  wire [6:0] _T_1983 = _T_509 ? 7'h70 : _T_1982; // @[Lookup.scala 33:37]
  wire [6:0] _T_1984 = _T_507 ? 7'h68 : _T_1983; // @[Lookup.scala 33:37]
  wire [6:0] _T_1985 = _T_505 ? 7'h60 : _T_1984; // @[Lookup.scala 33:37]
  wire [6:0] _T_1986 = _T_503 ? 7'h58 : _T_1985; // @[Lookup.scala 33:37]
  wire [6:0] _T_1987 = _T_501 ? 7'h78 : _T_1986; // @[Lookup.scala 33:37]
  wire [6:0] _T_1988 = _T_499 ? 7'h67 : _T_1987; // @[Lookup.scala 33:37]
  wire [6:0] _T_1989 = _T_497 ? 7'h3 : _T_1988; // @[Lookup.scala 33:37]
  wire [6:0] _T_1990 = _T_495 ? 7'h73 : _T_1989; // @[Lookup.scala 33:37]
  wire [6:0] _T_1991 = _T_493 ? 7'h12 : _T_1990; // @[Lookup.scala 33:37]
  wire [6:0] _T_1992 = _T_491 ? 7'h70 : _T_1991; // @[Lookup.scala 33:37]
  wire [6:0] _T_1993 = _T_489 ? 7'h19 : _T_1992; // @[Lookup.scala 33:37]
  wire [6:0] _T_1994 = _T_487 ? 7'h11 : _T_1993; // @[Lookup.scala 33:37]
  wire [6:0] _T_1995 = _T_485 ? 7'h18 : _T_1994; // @[Lookup.scala 33:37]
  wire [6:0] _T_1996 = _T_483 ? 7'h10 : _T_1995; // @[Lookup.scala 33:37]
  wire [6:0] _T_1997 = _T_481 ? 7'h13 : _T_1996; // @[Lookup.scala 33:37]
  wire [6:0] _T_1998 = _T_479 ? 7'h3f : _T_1997; // @[Lookup.scala 33:37]
  wire [6:0] _T_1999 = _T_477 ? 7'h37 : _T_1998; // @[Lookup.scala 33:37]
  wire [6:0] _T_2000 = _T_475 ? 7'h9 : _T_1999; // @[Lookup.scala 33:37]
  wire [6:0] _T_2001 = _T_473 ? 7'h1 : _T_2000; // @[Lookup.scala 33:37]
  wire [6:0] _T_2002 = _T_471 ? 7'h8 : _T_2001; // @[Lookup.scala 33:37]
  wire [6:0] _T_2003 = _T_469 ? 7'h0 : _T_2002; // @[Lookup.scala 33:37]
  wire [6:0] _T_2004 = _T_467 ? 7'hb : _T_2003; // @[Lookup.scala 33:37]
  wire [6:0] _T_2005 = _T_465 ? 7'h3 : _T_2004; // @[Lookup.scala 33:37]
  wire [6:0] _T_2006 = _T_463 ? 7'ha : _T_2005; // @[Lookup.scala 33:37]
  wire [6:0] _T_2007 = _T_461 ? 7'h2 : _T_2006; // @[Lookup.scala 33:37]
  wire [6:0] _T_2008 = _T_459 ? 7'h59 : _T_2007; // @[Lookup.scala 33:37]
  wire [6:0] _T_2009 = _T_457 ? 7'h51 : _T_2008; // @[Lookup.scala 33:37]
  wire [6:0] _T_2010 = _T_455 ? 7'h49 : _T_2009; // @[Lookup.scala 33:37]
  wire [6:0] _T_2011 = _T_453 ? 7'h41 : _T_2010; // @[Lookup.scala 33:37]
  wire [6:0] _T_2012 = _T_451 ? 7'h58 : _T_2011; // @[Lookup.scala 33:37]
  wire [6:0] _T_2013 = _T_449 ? 7'h50 : _T_2012; // @[Lookup.scala 33:37]
  wire [6:0] _T_2014 = _T_447 ? 7'h48 : _T_2013; // @[Lookup.scala 33:37]
  wire [6:0] _T_2015 = _T_445 ? 7'h40 : _T_2014; // @[Lookup.scala 33:37]
  wire [6:0] _T_2016 = _T_443 ? 7'h7f : _T_2015; // @[Lookup.scala 33:37]
  wire [6:0] _T_2017 = _T_441 ? 7'h7e : _T_2016; // @[Lookup.scala 33:37]
  wire [6:0] _T_2018 = _T_439 ? 7'h1f : _T_2017; // @[Lookup.scala 33:37]
  wire [6:0] _T_2019 = _T_437 ? 7'h17 : _T_2018; // @[Lookup.scala 33:37]
  wire [6:0] _T_2020 = _T_435 ? 7'hf : _T_2019; // @[Lookup.scala 33:37]
  wire [6:0] _T_2021 = _T_433 ? 7'h7 : _T_2020; // @[Lookup.scala 33:37]
  wire [6:0] _T_2022 = _T_431 ? 7'h4d : _T_2021; // @[Lookup.scala 33:37]
  wire [6:0] _T_2023 = _T_429 ? 7'h4c : _T_2022; // @[Lookup.scala 33:37]
  wire [6:0] _T_2024 = _T_427 ? 7'h45 : _T_2023; // @[Lookup.scala 33:37]
  wire [6:0] _T_2025 = _T_425 ? 7'h44 : _T_2024; // @[Lookup.scala 33:37]
  wire [6:0] _T_2026 = _T_423 ? 7'h49 : _T_2025; // @[Lookup.scala 33:37]
  wire [6:0] _T_2027 = _T_421 ? 7'h48 : _T_2026; // @[Lookup.scala 33:37]
  wire [6:0] _T_2028 = _T_419 ? 7'h41 : _T_2027; // @[Lookup.scala 33:37]
  wire [6:0] _T_2029 = _T_417 ? 7'h40 : _T_2028; // @[Lookup.scala 33:37]
  wire [6:0] _T_2030 = _T_415 ? 7'h1f : _T_2029; // @[Lookup.scala 33:37]
  wire [6:0] _T_2031 = _T_413 ? 7'h17 : _T_2030; // @[Lookup.scala 33:37]
  wire [6:0] _T_2032 = _T_411 ? 7'hf : _T_2031; // @[Lookup.scala 33:37]
  wire [6:0] _T_2033 = _T_409 ? 7'h7 : _T_2032; // @[Lookup.scala 33:37]
  wire [6:0] _T_2034 = _T_407 ? 7'h27 : _T_2033; // @[Lookup.scala 33:37]
  wire [6:0] _T_2035 = _T_405 ? 7'h1e : _T_2034; // @[Lookup.scala 33:37]
  wire [6:0] _T_2036 = _T_403 ? 7'h16 : _T_2035; // @[Lookup.scala 33:37]
  wire [6:0] _T_2037 = _T_401 ? 7'he : _T_2036; // @[Lookup.scala 33:37]
  wire [6:0] _T_2038 = _T_399 ? 7'h6 : _T_2037; // @[Lookup.scala 33:37]
  wire [6:0] _T_2039 = _T_397 ? 7'h26 : _T_2038; // @[Lookup.scala 33:37]
  wire [6:0] _T_2040 = _T_395 ? 7'h33 : _T_2039; // @[Lookup.scala 33:37]
  wire [6:0] _T_2041 = _T_393 ? 7'h2b : _T_2040; // @[Lookup.scala 33:37]
  wire [6:0] _T_2042 = _T_391 ? 7'h32 : _T_2041; // @[Lookup.scala 33:37]
  wire [6:0] _T_2043 = _T_389 ? 7'h2a : _T_2042; // @[Lookup.scala 33:37]
  wire [6:0] _T_2044 = _T_387 ? 7'h31 : _T_2043; // @[Lookup.scala 33:37]
  wire [6:0] _T_2045 = _T_385 ? 7'h29 : _T_2044; // @[Lookup.scala 33:37]
  wire [6:0] _T_2046 = _T_383 ? 7'h30 : _T_2045; // @[Lookup.scala 33:37]
  wire [6:0] _T_2047 = _T_381 ? 7'h28 : _T_2046; // @[Lookup.scala 33:37]
  wire [6:0] _T_2048 = _T_379 ? 7'h37 : _T_2047; // @[Lookup.scala 33:37]
  wire [6:0] _T_2049 = _T_377 ? 7'h2f : _T_2048; // @[Lookup.scala 33:37]
  wire [6:0] _T_2050 = _T_375 ? 7'h36 : _T_2049; // @[Lookup.scala 33:37]
  wire [6:0] _T_2051 = _T_373 ? 7'h2e : _T_2050; // @[Lookup.scala 33:37]
  wire [6:0] _T_2052 = _T_371 ? 7'h35 : _T_2051; // @[Lookup.scala 33:37]
  wire [6:0] _T_2053 = _T_369 ? 7'h2d : _T_2052; // @[Lookup.scala 33:37]
  wire [6:0] _T_2054 = _T_367 ? 7'h34 : _T_2053; // @[Lookup.scala 33:37]
  wire [6:0] _T_2055 = _T_365 ? 7'h2c : _T_2054; // @[Lookup.scala 33:37]
  wire [6:0] _T_2056 = _T_363 ? 7'h33 : _T_2055; // @[Lookup.scala 33:37]
  wire [6:0] _T_2057 = _T_361 ? 7'h2b : _T_2056; // @[Lookup.scala 33:37]
  wire [6:0] _T_2058 = _T_359 ? 7'h32 : _T_2057; // @[Lookup.scala 33:37]
  wire [6:0] _T_2059 = _T_357 ? 7'h2a : _T_2058; // @[Lookup.scala 33:37]
  wire [6:0] _T_2060 = _T_355 ? 7'h31 : _T_2059; // @[Lookup.scala 33:37]
  wire [6:0] _T_2061 = _T_353 ? 7'h29 : _T_2060; // @[Lookup.scala 33:37]
  wire [6:0] _T_2062 = _T_351 ? 7'h30 : _T_2061; // @[Lookup.scala 33:37]
  wire [6:0] _T_2063 = _T_349 ? 7'h28 : _T_2062; // @[Lookup.scala 33:37]
  wire [6:0] _T_2064 = _T_347 ? 7'h1b : _T_2063; // @[Lookup.scala 33:37]
  wire [6:0] _T_2065 = _T_345 ? 7'h13 : _T_2064; // @[Lookup.scala 33:37]
  wire [6:0] _T_2066 = _T_343 ? 7'hb : _T_2065; // @[Lookup.scala 33:37]
  wire [6:0] _T_2067 = _T_341 ? 7'h3 : _T_2066; // @[Lookup.scala 33:37]
  wire [6:0] _T_2068 = _T_339 ? 7'h23 : _T_2067; // @[Lookup.scala 33:37]
  wire [6:0] _T_2069 = _T_337 ? 7'h1a : _T_2068; // @[Lookup.scala 33:37]
  wire [6:0] _T_2070 = _T_335 ? 7'h12 : _T_2069; // @[Lookup.scala 33:37]
  wire [6:0] _T_2071 = _T_333 ? 7'ha : _T_2070; // @[Lookup.scala 33:37]
  wire [6:0] _T_2072 = _T_331 ? 7'h2 : _T_2071; // @[Lookup.scala 33:37]
  wire [6:0] _T_2073 = _T_329 ? 7'h22 : _T_2072; // @[Lookup.scala 33:37]
  wire [6:0] _T_2074 = _T_327 ? 7'h19 : _T_2073; // @[Lookup.scala 33:37]
  wire [6:0] _T_2075 = _T_325 ? 7'h11 : _T_2074; // @[Lookup.scala 33:37]
  wire [6:0] _T_2076 = _T_323 ? 7'h9 : _T_2075; // @[Lookup.scala 33:37]
  wire [6:0] _T_2077 = _T_321 ? 7'h1 : _T_2076; // @[Lookup.scala 33:37]
  wire [6:0] _T_2078 = _T_319 ? 7'h21 : _T_2077; // @[Lookup.scala 33:37]
  wire [6:0] _T_2079 = _T_317 ? 7'h18 : _T_2078; // @[Lookup.scala 33:37]
  wire [6:0] _T_2080 = _T_315 ? 7'h10 : _T_2079; // @[Lookup.scala 33:37]
  wire [6:0] _T_2081 = _T_313 ? 7'h8 : _T_2080; // @[Lookup.scala 33:37]
  wire [6:0] _T_2082 = _T_311 ? 7'h0 : _T_2081; // @[Lookup.scala 33:37]
  wire [6:0] _T_2083 = _T_309 ? 7'h20 : _T_2082; // @[Lookup.scala 33:37]
  wire [6:0] _T_2084 = _T_307 ? 7'h1b : _T_2083; // @[Lookup.scala 33:37]
  wire [6:0] _T_2085 = _T_305 ? 7'h13 : _T_2084; // @[Lookup.scala 33:37]
  wire [6:0] _T_2086 = _T_303 ? 7'hb : _T_2085; // @[Lookup.scala 33:37]
  wire [6:0] _T_2087 = _T_301 ? 7'h3 : _T_2086; // @[Lookup.scala 33:37]
  wire [6:0] _T_2088 = _T_299 ? 7'h23 : _T_2087; // @[Lookup.scala 33:37]
  wire [6:0] _T_2089 = _T_297 ? 7'h1a : _T_2088; // @[Lookup.scala 33:37]
  wire [6:0] _T_2090 = _T_295 ? 7'h12 : _T_2089; // @[Lookup.scala 33:37]
  wire [6:0] _T_2091 = _T_293 ? 7'ha : _T_2090; // @[Lookup.scala 33:37]
  wire [6:0] _T_2092 = _T_291 ? 7'h2 : _T_2091; // @[Lookup.scala 33:37]
  wire [6:0] _T_2093 = _T_289 ? 7'h22 : _T_2092; // @[Lookup.scala 33:37]
  wire [6:0] _T_2094 = _T_287 ? 7'h1d : _T_2093; // @[Lookup.scala 33:37]
  wire [6:0] _T_2095 = _T_285 ? 7'h15 : _T_2094; // @[Lookup.scala 33:37]
  wire [6:0] _T_2096 = _T_283 ? 7'hd : _T_2095; // @[Lookup.scala 33:37]
  wire [6:0] _T_2097 = _T_281 ? 7'h5 : _T_2096; // @[Lookup.scala 33:37]
  wire [6:0] _T_2098 = _T_279 ? 7'h25 : _T_2097; // @[Lookup.scala 33:37]
  wire [6:0] _T_2099 = _T_277 ? 7'h1c : _T_2098; // @[Lookup.scala 33:37]
  wire [6:0] _T_2100 = _T_275 ? 7'h14 : _T_2099; // @[Lookup.scala 33:37]
  wire [6:0] _T_2101 = _T_273 ? 7'hc : _T_2100; // @[Lookup.scala 33:37]
  wire [6:0] _T_2102 = _T_271 ? 7'h4 : _T_2101; // @[Lookup.scala 33:37]
  wire [6:0] _T_2103 = _T_269 ? 7'h24 : _T_2102; // @[Lookup.scala 33:37]
  wire [6:0] _T_2104 = _T_267 ? 7'h19 : _T_2103; // @[Lookup.scala 33:37]
  wire [6:0] _T_2105 = _T_265 ? 7'h11 : _T_2104; // @[Lookup.scala 33:37]
  wire [6:0] _T_2106 = _T_263 ? 7'h9 : _T_2105; // @[Lookup.scala 33:37]
  wire [6:0] _T_2107 = _T_261 ? 7'h1 : _T_2106; // @[Lookup.scala 33:37]
  wire [6:0] _T_2108 = _T_259 ? 7'h21 : _T_2107; // @[Lookup.scala 33:37]
  wire [6:0] _T_2109 = _T_257 ? 7'h18 : _T_2108; // @[Lookup.scala 33:37]
  wire [6:0] _T_2110 = _T_255 ? 7'h10 : _T_2109; // @[Lookup.scala 33:37]
  wire [6:0] _T_2111 = _T_253 ? 7'h8 : _T_2110; // @[Lookup.scala 33:37]
  wire [6:0] _T_2112 = _T_251 ? 7'h0 : _T_2111; // @[Lookup.scala 33:37]
  wire [6:0] _T_2113 = _T_249 ? 7'h20 : _T_2112; // @[Lookup.scala 33:37]
  wire [6:0] _T_2114 = _T_247 ? 7'h1 : _T_2113; // @[Lookup.scala 33:37]
  wire [6:0] _T_2115 = _T_245 ? 7'h7 : _T_2114; // @[Lookup.scala 33:37]
  wire [6:0] _T_2116 = _T_243 ? 7'h6 : _T_2115; // @[Lookup.scala 33:37]
  wire [6:0] _T_2117 = _T_241 ? 7'h5 : _T_2116; // @[Lookup.scala 33:37]
  wire [6:0] _T_2118 = _T_239 ? 7'h3 : _T_2117; // @[Lookup.scala 33:37]
  wire [6:0] _T_2119 = _T_237 ? 7'h2 : _T_2118; // @[Lookup.scala 33:37]
  wire [6:0] _T_2120 = _T_235 ? 7'h1 : _T_2119; // @[Lookup.scala 33:37]
  wire [6:0] _T_2121 = _T_233 ? 7'h32 : _T_2120; // @[Lookup.scala 33:37]
  wire [6:0] _T_2122 = _T_231 ? 7'h31 : _T_2121; // @[Lookup.scala 33:37]
  wire [6:0] _T_2123 = _T_229 ? 7'h30 : _T_2122; // @[Lookup.scala 33:37]
  wire [6:0] _T_2124 = _T_227 ? 7'h37 : _T_2123; // @[Lookup.scala 33:37]
  wire [6:0] _T_2125 = _T_225 ? 7'h26 : _T_2124; // @[Lookup.scala 33:37]
  wire [6:0] _T_2126 = _T_223 ? 7'h25 : _T_2125; // @[Lookup.scala 33:37]
  wire [6:0] _T_2127 = _T_221 ? 7'h24 : _T_2126; // @[Lookup.scala 33:37]
  wire [6:0] _T_2128 = _T_219 ? 7'h63 : _T_2127; // @[Lookup.scala 33:37]
  wire [6:0] _T_2129 = _T_217 ? 7'h22 : _T_2128; // @[Lookup.scala 33:37]
  wire [6:0] _T_2130 = _T_215 ? 7'h21 : _T_2129; // @[Lookup.scala 33:37]
  wire [6:0] _T_2131 = _T_213 ? 7'h21 : _T_2130; // @[Lookup.scala 33:37]
  wire [6:0] _T_2132 = _T_211 ? 7'h20 : _T_2131; // @[Lookup.scala 33:37]
  wire [6:0] _T_2133 = _T_209 ? 7'h20 : _T_2132; // @[Lookup.scala 33:37]
  wire [6:0] _T_2134 = _T_207 ? 7'h2 : _T_2133; // @[Lookup.scala 33:37]
  wire [6:0] _T_2135 = _T_205 ? 7'h0 : _T_2134; // @[Lookup.scala 33:37]
  wire [6:0] _T_2136 = _T_203 ? 7'h40 : _T_2135; // @[Lookup.scala 33:37]
  wire [6:0] _T_2137 = _T_201 ? 7'h0 : _T_2136; // @[Lookup.scala 33:37]
  wire [6:0] _T_2138 = _T_199 ? 7'h0 : _T_2137; // @[Lookup.scala 33:37]
  wire [6:0] _T_2139 = _T_197 ? 7'h0 : _T_2138; // @[Lookup.scala 33:37]
  wire [6:0] _T_2140 = _T_195 ? 7'h0 : _T_2139; // @[Lookup.scala 33:37]
  wire [6:0] _T_2141 = _T_193 ? 7'hb : _T_2140; // @[Lookup.scala 33:37]
  wire [6:0] _T_2142 = _T_191 ? 7'ha : _T_2141; // @[Lookup.scala 33:37]
  wire [6:0] _T_2143 = _T_189 ? 7'h40 : _T_2142; // @[Lookup.scala 33:37]
  wire [6:0] _T_2144 = _T_187 ? 7'h5a : _T_2143; // @[Lookup.scala 33:37]
  wire [6:0] _T_2145 = _T_185 ? 7'h0 : _T_2144; // @[Lookup.scala 33:37]
  wire [6:0] _T_2146 = _T_183 ? 7'h40 : _T_2145; // @[Lookup.scala 33:37]
  wire [6:0] _T_2147 = _T_181 ? 7'h5a : _T_2146; // @[Lookup.scala 33:37]
  wire [6:0] _T_2148 = _T_179 ? 7'h3 : _T_2147; // @[Lookup.scala 33:37]
  wire [6:0] _T_2149 = _T_177 ? 7'h2 : _T_2148; // @[Lookup.scala 33:37]
  wire [6:0] _T_2150 = _T_175 ? 7'h1 : _T_2149; // @[Lookup.scala 33:37]
  wire [6:0] _T_2151 = _T_173 ? 7'h11 : _T_2150; // @[Lookup.scala 33:37]
  wire [6:0] _T_2152 = _T_171 ? 7'h10 : _T_2151; // @[Lookup.scala 33:37]
  wire [6:0] _T_2153 = _T_169 ? 7'h58 : _T_2152; // @[Lookup.scala 33:37]
  wire [6:0] _T_2154 = _T_167 ? 7'h60 : _T_2153; // @[Lookup.scala 33:37]
  wire [6:0] _T_2155 = _T_165 ? 7'h28 : _T_2154; // @[Lookup.scala 33:37]
  wire [6:0] _T_2156 = _T_163 ? 7'h7 : _T_2155; // @[Lookup.scala 33:37]
  wire [6:0] _T_2157 = _T_161 ? 7'h6 : _T_2156; // @[Lookup.scala 33:37]
  wire [6:0] _T_2158 = _T_159 ? 7'h4 : _T_2157; // @[Lookup.scala 33:37]
  wire [6:0] _T_2159 = _T_157 ? 7'h8 : _T_2158; // @[Lookup.scala 33:37]
  wire [6:0] _T_2160 = _T_155 ? 7'h7 : _T_2159; // @[Lookup.scala 33:37]
  wire [6:0] _T_2161 = _T_153 ? 7'hd : _T_2160; // @[Lookup.scala 33:37]
  wire [6:0] _T_2162 = _T_151 ? 7'h5 : _T_2161; // @[Lookup.scala 33:37]
  wire [6:0] _T_2163 = _T_149 ? 7'h40 : _T_2162; // @[Lookup.scala 33:37]
  wire [6:0] _T_2164 = _T_147 ? 7'h40 : _T_2163; // @[Lookup.scala 33:37]
  wire [6:0] _T_2165 = _T_145 ? 7'h40 : _T_2164; // @[Lookup.scala 33:37]
  wire [6:0] _T_2166 = _T_143 ? 7'h60 : _T_2165; // @[Lookup.scala 33:37]
  wire [6:0] _T_2167 = _T_141 ? 7'h40 : _T_2166; // @[Lookup.scala 33:37]
  wire [6:0] _T_2168 = _T_139 ? 7'h40 : _T_2167; // @[Lookup.scala 33:37]
  wire [6:0] _T_2169 = _T_137 ? 7'hb : _T_2168; // @[Lookup.scala 33:37]
  wire [6:0] _T_2170 = _T_135 ? 7'ha : _T_2169; // @[Lookup.scala 33:37]
  wire [6:0] _T_2171 = _T_133 ? 7'h3 : _T_2170; // @[Lookup.scala 33:37]
  wire [6:0] _T_2172 = _T_131 ? 7'h2 : _T_2171; // @[Lookup.scala 33:37]
  wire [6:0] _T_2173 = _T_129 ? 7'h40 : _T_2172; // @[Lookup.scala 33:37]
  wire [6:0] _T_2174 = _T_127 ? 7'h0 : _T_2173; // @[Lookup.scala 33:37]
  wire [6:0] _T_2175 = _T_125 ? 7'hf : _T_2174; // @[Lookup.scala 33:37]
  wire [6:0] _T_2176 = _T_123 ? 7'he : _T_2175; // @[Lookup.scala 33:37]
  wire [6:0] _T_2177 = _T_121 ? 7'hd : _T_2176; // @[Lookup.scala 33:37]
  wire [6:0] _T_2178 = _T_119 ? 7'hc : _T_2177; // @[Lookup.scala 33:37]
  wire [6:0] _T_2179 = _T_117 ? 7'h8 : _T_2178; // @[Lookup.scala 33:37]
  wire [6:0] _T_2180 = _T_115 ? 7'h7 : _T_2179; // @[Lookup.scala 33:37]
  wire [6:0] _T_2181 = _T_113 ? 7'h6 : _T_2180; // @[Lookup.scala 33:37]
  wire [6:0] _T_2182 = _T_111 ? 7'h5 : _T_2181; // @[Lookup.scala 33:37]
  wire [6:0] _T_2183 = _T_109 ? 7'h4 : _T_2182; // @[Lookup.scala 33:37]
  wire [6:0] _T_2184 = _T_107 ? 7'h3 : _T_2183; // @[Lookup.scala 33:37]
  wire [6:0] _T_2185 = _T_105 ? 7'h2 : _T_2184; // @[Lookup.scala 33:37]
  wire [6:0] _T_2186 = _T_103 ? 7'h1 : _T_2185; // @[Lookup.scala 33:37]
  wire [6:0] _T_2187 = _T_101 ? 7'h0 : _T_2186; // @[Lookup.scala 33:37]
  wire [6:0] _T_2188 = _T_99 ? 7'h2 : _T_2187; // @[Lookup.scala 33:37]
  wire [6:0] _T_2189 = _T_97 ? 7'hb : _T_2188; // @[Lookup.scala 33:37]
  wire [6:0] _T_2190 = _T_95 ? 7'h3 : _T_2189; // @[Lookup.scala 33:37]
  wire [6:0] _T_2191 = _T_93 ? 7'h6 : _T_2190; // @[Lookup.scala 33:37]
  wire [6:0] _T_2192 = _T_91 ? 7'h28 : _T_2191; // @[Lookup.scala 33:37]
  wire [6:0] _T_2193 = _T_89 ? 7'h60 : _T_2192; // @[Lookup.scala 33:37]
  wire [6:0] _T_2194 = _T_87 ? 7'h2d : _T_2193; // @[Lookup.scala 33:37]
  wire [6:0] _T_2195 = _T_85 ? 7'h25 : _T_2194; // @[Lookup.scala 33:37]
  wire [6:0] _T_2196 = _T_83 ? 7'h21 : _T_2195; // @[Lookup.scala 33:37]
  wire [6:0] _T_2197 = _T_81 ? 7'h2d : _T_2196; // @[Lookup.scala 33:37]
  wire [6:0] _T_2198 = _T_79 ? 7'h25 : _T_2197; // @[Lookup.scala 33:37]
  wire [6:0] _T_2199 = _T_77 ? 7'h21 : _T_2198; // @[Lookup.scala 33:37]
  wire [6:0] _T_2200 = _T_75 ? 7'h60 : _T_2199; // @[Lookup.scala 33:37]
  wire [6:0] _T_2201 = _T_73 ? 7'ha : _T_2200; // @[Lookup.scala 33:37]
  wire [6:0] _T_2202 = _T_71 ? 7'h9 : _T_2201; // @[Lookup.scala 33:37]
  wire [6:0] _T_2203 = _T_69 ? 7'h8 : _T_2202; // @[Lookup.scala 33:37]
  wire [6:0] _T_2204 = _T_67 ? 7'h5 : _T_2203; // @[Lookup.scala 33:37]
  wire [6:0] _T_2205 = _T_65 ? 7'h4 : _T_2204; // @[Lookup.scala 33:37]
  wire [6:0] _T_2206 = _T_63 ? 7'h2 : _T_2205; // @[Lookup.scala 33:37]
  wire [6:0] _T_2207 = _T_61 ? 7'h1 : _T_2206; // @[Lookup.scala 33:37]
  wire [6:0] _T_2208 = _T_59 ? 7'h0 : _T_2207; // @[Lookup.scala 33:37]
  wire [6:0] _T_2209 = _T_57 ? 7'h17 : _T_2208; // @[Lookup.scala 33:37]
  wire [6:0] _T_2210 = _T_55 ? 7'h16 : _T_2209; // @[Lookup.scala 33:37]
  wire [6:0] _T_2211 = _T_53 ? 7'h15 : _T_2210; // @[Lookup.scala 33:37]
  wire [6:0] _T_2212 = _T_51 ? 7'h14 : _T_2211; // @[Lookup.scala 33:37]
  wire [6:0] _T_2213 = _T_49 ? 7'h11 : _T_2212; // @[Lookup.scala 33:37]
  wire [6:0] _T_2214 = _T_47 ? 7'h10 : _T_2213; // @[Lookup.scala 33:37]
  wire [6:0] _T_2215 = _T_45 ? 7'h5a : _T_2214; // @[Lookup.scala 33:37]
  wire [6:0] _T_2216 = _T_43 ? 7'h58 : _T_2215; // @[Lookup.scala 33:37]
  wire [6:0] _T_2217 = _T_41 ? 7'h40 : _T_2216; // @[Lookup.scala 33:37]
  wire [6:0] _T_2218 = _T_39 ? 7'h40 : _T_2217; // @[Lookup.scala 33:37]
  wire [6:0] _T_2219 = _T_37 ? 7'hd : _T_2218; // @[Lookup.scala 33:37]
  wire [6:0] _T_2220 = _T_35 ? 7'h8 : _T_2219; // @[Lookup.scala 33:37]
  wire [6:0] _T_2221 = _T_33 ? 7'h7 : _T_2220; // @[Lookup.scala 33:37]
  wire [6:0] _T_2222 = _T_31 ? 7'h6 : _T_2221; // @[Lookup.scala 33:37]
  wire [6:0] _T_2223 = _T_29 ? 7'h5 : _T_2222; // @[Lookup.scala 33:37]
  wire [6:0] _T_2224 = _T_27 ? 7'h4 : _T_2223; // @[Lookup.scala 33:37]
  wire [6:0] _T_2225 = _T_25 ? 7'h3 : _T_2224; // @[Lookup.scala 33:37]
  wire [6:0] _T_2226 = _T_23 ? 7'h2 : _T_2225; // @[Lookup.scala 33:37]
  wire [6:0] _T_2227 = _T_21 ? 7'h1 : _T_2226; // @[Lookup.scala 33:37]
  wire [6:0] _T_2228 = _T_19 ? 7'h40 : _T_2227; // @[Lookup.scala 33:37]
  wire [6:0] _T_2229 = _T_17 ? 7'hd : _T_2228; // @[Lookup.scala 33:37]
  wire [6:0] _T_2230 = _T_15 ? 7'h7 : _T_2229; // @[Lookup.scala 33:37]
  wire [6:0] _T_2231 = _T_13 ? 7'h6 : _T_2230; // @[Lookup.scala 33:37]
  wire [6:0] _T_2232 = _T_11 ? 7'h5 : _T_2231; // @[Lookup.scala 33:37]
  wire [6:0] _T_2233 = _T_9 ? 7'h4 : _T_2232; // @[Lookup.scala 33:37]
  wire [6:0] _T_2234 = _T_7 ? 7'h3 : _T_2233; // @[Lookup.scala 33:37]
  wire [6:0] _T_2235 = _T_5 ? 7'h2 : _T_2234; // @[Lookup.scala 33:37]
  wire [6:0] _T_2236 = _T_3 ? 7'h1 : _T_2235; // @[Lookup.scala 33:37]
  wire [6:0] decodeList_2 = _T_1 ? 7'h40 : _T_2236; // @[Lookup.scala 33:37]
  wire [11:0] intrVec = intrVecIDU[11:0];
  wire  hasIntr = |intrVec; // @[IDU.scala 191:22]
  wire [4:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 5'h0 : decodeList_0; // @[IDU.scala 38:75]
  wire [3:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h1 : decodeList_1; // @[IDU.scala 38:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[IDU.scala 38:75]
  wire  isRVC = io_in_bits_instr[1:0] != 2'h3; // @[IDU.scala 40:45]
  wire [4:0] _T_2310 = _T_193 ? 5'h3 : 5'h10; // @[Lookup.scala 33:37]
  wire [4:0] _T_2311 = _T_191 ? 5'h2 : _T_2310; // @[Lookup.scala 33:37]
  wire [4:0] _T_2312 = _T_189 ? 5'h10 : _T_2311; // @[Lookup.scala 33:37]
  wire [4:0] _T_2313 = _T_187 ? 5'h10 : _T_2312; // @[Lookup.scala 33:37]
  wire [4:0] _T_2314 = _T_185 ? 5'hf : _T_2313; // @[Lookup.scala 33:37]
  wire [4:0] _T_2315 = _T_183 ? 5'h10 : _T_2314; // @[Lookup.scala 33:37]
  wire [4:0] _T_2316 = _T_181 ? 5'h10 : _T_2315; // @[Lookup.scala 33:37]
  wire [4:0] _T_2317 = _T_179 ? 5'h1 : _T_2316; // @[Lookup.scala 33:37]
  wire [4:0] _T_2318 = _T_177 ? 5'h0 : _T_2317; // @[Lookup.scala 33:37]
  wire [4:0] _T_2319 = _T_175 ? 5'ha : _T_2318; // @[Lookup.scala 33:37]
  wire [4:0] _T_2320 = _T_173 ? 5'h9 : _T_2319; // @[Lookup.scala 33:37]
  wire [4:0] _T_2321 = _T_171 ? 5'h9 : _T_2320; // @[Lookup.scala 33:37]
  wire [4:0] _T_2322 = _T_169 ? 5'h8 : _T_2321; // @[Lookup.scala 33:37]
  wire [4:0] _T_2323 = _T_167 ? 5'h10 : _T_2322; // @[Lookup.scala 33:37]
  wire [4:0] _T_2324 = _T_165 ? 5'h10 : _T_2323; // @[Lookup.scala 33:37]
  wire [4:0] _T_2325 = _T_163 ? 5'h10 : _T_2324; // @[Lookup.scala 33:37]
  wire [4:0] _T_2326 = _T_161 ? 5'h10 : _T_2325; // @[Lookup.scala 33:37]
  wire [4:0] _T_2327 = _T_159 ? 5'h10 : _T_2326; // @[Lookup.scala 33:37]
  wire [4:0] _T_2328 = _T_157 ? 5'h10 : _T_2327; // @[Lookup.scala 33:37]
  wire [4:0] _T_2329 = _T_155 ? 5'ha : _T_2328; // @[Lookup.scala 33:37]
  wire [4:0] _T_2330 = _T_153 ? 5'ha : _T_2329; // @[Lookup.scala 33:37]
  wire [4:0] _T_2331 = _T_151 ? 5'ha : _T_2330; // @[Lookup.scala 33:37]
  wire [4:0] _T_2332 = _T_149 ? 5'hb : _T_2331; // @[Lookup.scala 33:37]
  wire [4:0] _T_2333 = _T_147 ? 5'hd : _T_2332; // @[Lookup.scala 33:37]
  wire [4:0] _T_2334 = _T_145 ? 5'ha : _T_2333; // @[Lookup.scala 33:37]
  wire [4:0] _T_2335 = _T_143 ? 5'hc : _T_2334; // @[Lookup.scala 33:37]
  wire [4:0] _T_2336 = _T_141 ? 5'hc : _T_2335; // @[Lookup.scala 33:37]
  wire [4:0] _T_2337 = _T_139 ? 5'h10 : _T_2336; // @[Lookup.scala 33:37]
  wire [4:0] _T_2338 = _T_137 ? 5'h5 : _T_2337; // @[Lookup.scala 33:37]
  wire [4:0] _T_2339 = _T_135 ? 5'h4 : _T_2338; // @[Lookup.scala 33:37]
  wire [4:0] _T_2340 = _T_133 ? 5'h7 : _T_2339; // @[Lookup.scala 33:37]
  wire [4:0] _T_2341 = _T_131 ? 5'h6 : _T_2340; // @[Lookup.scala 33:37]
  wire [4:0] rvcImmType = _T_129 ? 5'he : _T_2341; // @[Lookup.scala 33:37]
  wire [3:0] _T_2342 = _T_193 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_2343 = _T_191 ? 4'h9 : _T_2342; // @[Lookup.scala 33:37]
  wire [3:0] _T_2344 = _T_189 ? 4'h2 : _T_2343; // @[Lookup.scala 33:37]
  wire [3:0] _T_2345 = _T_187 ? 4'h4 : _T_2344; // @[Lookup.scala 33:37]
  wire [3:0] _T_2346 = _T_185 ? 4'h0 : _T_2345; // @[Lookup.scala 33:37]
  wire [3:0] _T_2347 = _T_183 ? 4'h5 : _T_2346; // @[Lookup.scala 33:37]
  wire [3:0] _T_2348 = _T_181 ? 4'h4 : _T_2347; // @[Lookup.scala 33:37]
  wire [3:0] _T_2349 = _T_179 ? 4'h9 : _T_2348; // @[Lookup.scala 33:37]
  wire [3:0] _T_2350 = _T_177 ? 4'h9 : _T_2349; // @[Lookup.scala 33:37]
  wire [3:0] _T_2351 = _T_175 ? 4'h2 : _T_2350; // @[Lookup.scala 33:37]
  wire [3:0] _T_2352 = _T_173 ? 4'h6 : _T_2351; // @[Lookup.scala 33:37]
  wire [3:0] _T_2353 = _T_171 ? 4'h6 : _T_2352; // @[Lookup.scala 33:37]
  wire [3:0] _T_2354 = _T_169 ? 4'h0 : _T_2353; // @[Lookup.scala 33:37]
  wire [3:0] _T_2355 = _T_167 ? 4'h6 : _T_2354; // @[Lookup.scala 33:37]
  wire [3:0] _T_2356 = _T_165 ? 4'h6 : _T_2355; // @[Lookup.scala 33:37]
  wire [3:0] _T_2357 = _T_163 ? 4'h6 : _T_2356; // @[Lookup.scala 33:37]
  wire [3:0] _T_2358 = _T_161 ? 4'h6 : _T_2357; // @[Lookup.scala 33:37]
  wire [3:0] _T_2359 = _T_159 ? 4'h6 : _T_2358; // @[Lookup.scala 33:37]
  wire [3:0] _T_2360 = _T_157 ? 4'h6 : _T_2359; // @[Lookup.scala 33:37]
  wire [3:0] _T_2361 = _T_155 ? 4'h6 : _T_2360; // @[Lookup.scala 33:37]
  wire [3:0] _T_2362 = _T_153 ? 4'h6 : _T_2361; // @[Lookup.scala 33:37]
  wire [3:0] _T_2363 = _T_151 ? 4'h6 : _T_2362; // @[Lookup.scala 33:37]
  wire [3:0] _T_2364 = _T_149 ? 4'h0 : _T_2363; // @[Lookup.scala 33:37]
  wire [3:0] _T_2365 = _T_147 ? 4'h9 : _T_2364; // @[Lookup.scala 33:37]
  wire [3:0] _T_2366 = _T_145 ? 4'h0 : _T_2365; // @[Lookup.scala 33:37]
  wire [3:0] _T_2367 = _T_143 ? 4'h2 : _T_2366; // @[Lookup.scala 33:37]
  wire [3:0] _T_2368 = _T_141 ? 4'h2 : _T_2367; // @[Lookup.scala 33:37]
  wire [3:0] _T_2369 = _T_139 ? 4'h0 : _T_2368; // @[Lookup.scala 33:37]
  wire [3:0] _T_2370 = _T_137 ? 4'h6 : _T_2369; // @[Lookup.scala 33:37]
  wire [3:0] _T_2371 = _T_135 ? 4'h6 : _T_2370; // @[Lookup.scala 33:37]
  wire [3:0] _T_2372 = _T_133 ? 4'h6 : _T_2371; // @[Lookup.scala 33:37]
  wire [3:0] _T_2373 = _T_131 ? 4'h6 : _T_2372; // @[Lookup.scala 33:37]
  wire [3:0] rvcSrc1Type = _T_129 ? 4'h9 : _T_2373; // @[Lookup.scala 33:37]
  wire [2:0] _T_2374 = _T_193 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_2375 = _T_191 ? 3'h5 : _T_2374; // @[Lookup.scala 33:37]
  wire [2:0] _T_2376 = _T_189 ? 3'h5 : _T_2375; // @[Lookup.scala 33:37]
  wire [2:0] _T_2377 = _T_187 ? 3'h0 : _T_2376; // @[Lookup.scala 33:37]
  wire [2:0] _T_2378 = _T_185 ? 3'h0 : _T_2377; // @[Lookup.scala 33:37]
  wire [2:0] _T_2379 = _T_183 ? 3'h0 : _T_2378; // @[Lookup.scala 33:37]
  wire [2:0] _T_2380 = _T_181 ? 3'h0 : _T_2379; // @[Lookup.scala 33:37]
  wire [2:0] _T_2381 = _T_179 ? 3'h0 : _T_2380; // @[Lookup.scala 33:37]
  wire [2:0] _T_2382 = _T_177 ? 3'h0 : _T_2381; // @[Lookup.scala 33:37]
  wire [2:0] _T_2383 = _T_175 ? 3'h0 : _T_2382; // @[Lookup.scala 33:37]
  wire [2:0] _T_2384 = _T_173 ? 3'h0 : _T_2383; // @[Lookup.scala 33:37]
  wire [2:0] _T_2385 = _T_171 ? 3'h0 : _T_2384; // @[Lookup.scala 33:37]
  wire [2:0] _T_2386 = _T_169 ? 3'h0 : _T_2385; // @[Lookup.scala 33:37]
  wire [2:0] _T_2387 = _T_167 ? 3'h7 : _T_2386; // @[Lookup.scala 33:37]
  wire [2:0] _T_2388 = _T_165 ? 3'h7 : _T_2387; // @[Lookup.scala 33:37]
  wire [2:0] _T_2389 = _T_163 ? 3'h7 : _T_2388; // @[Lookup.scala 33:37]
  wire [2:0] _T_2390 = _T_161 ? 3'h7 : _T_2389; // @[Lookup.scala 33:37]
  wire [2:0] _T_2391 = _T_159 ? 3'h7 : _T_2390; // @[Lookup.scala 33:37]
  wire [2:0] _T_2392 = _T_157 ? 3'h7 : _T_2391; // @[Lookup.scala 33:37]
  wire [2:0] _T_2393 = _T_155 ? 3'h0 : _T_2392; // @[Lookup.scala 33:37]
  wire [2:0] _T_2394 = _T_153 ? 3'h0 : _T_2393; // @[Lookup.scala 33:37]
  wire [2:0] _T_2395 = _T_151 ? 3'h0 : _T_2394; // @[Lookup.scala 33:37]
  wire [2:0] _T_2396 = _T_149 ? 3'h0 : _T_2395; // @[Lookup.scala 33:37]
  wire [2:0] _T_2397 = _T_147 ? 3'h0 : _T_2396; // @[Lookup.scala 33:37]
  wire [2:0] _T_2398 = _T_145 ? 3'h0 : _T_2397; // @[Lookup.scala 33:37]
  wire [2:0] _T_2399 = _T_143 ? 3'h0 : _T_2398; // @[Lookup.scala 33:37]
  wire [2:0] _T_2400 = _T_141 ? 3'h0 : _T_2399; // @[Lookup.scala 33:37]
  wire [2:0] _T_2401 = _T_139 ? 3'h0 : _T_2400; // @[Lookup.scala 33:37]
  wire [2:0] _T_2402 = _T_137 ? 3'h7 : _T_2401; // @[Lookup.scala 33:37]
  wire [2:0] _T_2403 = _T_135 ? 3'h7 : _T_2402; // @[Lookup.scala 33:37]
  wire [2:0] _T_2404 = _T_133 ? 3'h0 : _T_2403; // @[Lookup.scala 33:37]
  wire [2:0] _T_2405 = _T_131 ? 3'h0 : _T_2404; // @[Lookup.scala 33:37]
  wire [2:0] rvcSrc2Type = _T_129 ? 3'h0 : _T_2405; // @[Lookup.scala 33:37]
  wire [1:0] _T_2408 = _T_189 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_2409 = _T_187 ? 4'h8 : {{2'd0}, _T_2408}; // @[Lookup.scala 33:37]
  wire [3:0] _T_2410 = _T_185 ? 4'h0 : _T_2409; // @[Lookup.scala 33:37]
  wire [3:0] _T_2411 = _T_183 ? 4'h2 : _T_2410; // @[Lookup.scala 33:37]
  wire [3:0] _T_2412 = _T_181 ? 4'h0 : _T_2411; // @[Lookup.scala 33:37]
  wire [3:0] _T_2413 = _T_179 ? 4'h2 : _T_2412; // @[Lookup.scala 33:37]
  wire [3:0] _T_2414 = _T_177 ? 4'h2 : _T_2413; // @[Lookup.scala 33:37]
  wire [3:0] _T_2415 = _T_175 ? 4'h2 : _T_2414; // @[Lookup.scala 33:37]
  wire [3:0] _T_2416 = _T_173 ? 4'h0 : _T_2415; // @[Lookup.scala 33:37]
  wire [3:0] _T_2417 = _T_171 ? 4'h0 : _T_2416; // @[Lookup.scala 33:37]
  wire [3:0] _T_2418 = _T_169 ? 4'h0 : _T_2417; // @[Lookup.scala 33:37]
  wire [3:0] _T_2419 = _T_167 ? 4'h6 : _T_2418; // @[Lookup.scala 33:37]
  wire [3:0] _T_2420 = _T_165 ? 4'h6 : _T_2419; // @[Lookup.scala 33:37]
  wire [3:0] _T_2421 = _T_163 ? 4'h6 : _T_2420; // @[Lookup.scala 33:37]
  wire [3:0] _T_2422 = _T_161 ? 4'h6 : _T_2421; // @[Lookup.scala 33:37]
  wire [3:0] _T_2423 = _T_159 ? 4'h6 : _T_2422; // @[Lookup.scala 33:37]
  wire [3:0] _T_2424 = _T_157 ? 4'h6 : _T_2423; // @[Lookup.scala 33:37]
  wire [3:0] _T_2425 = _T_155 ? 4'h6 : _T_2424; // @[Lookup.scala 33:37]
  wire [3:0] _T_2426 = _T_153 ? 4'h6 : _T_2425; // @[Lookup.scala 33:37]
  wire [3:0] _T_2427 = _T_151 ? 4'h6 : _T_2426; // @[Lookup.scala 33:37]
  wire [3:0] _T_2428 = _T_149 ? 4'h2 : _T_2427; // @[Lookup.scala 33:37]
  wire [3:0] _T_2429 = _T_147 ? 4'h9 : _T_2428; // @[Lookup.scala 33:37]
  wire [3:0] _T_2430 = _T_145 ? 4'h2 : _T_2429; // @[Lookup.scala 33:37]
  wire [3:0] _T_2431 = _T_143 ? 4'h2 : _T_2430; // @[Lookup.scala 33:37]
  wire [3:0] _T_2432 = _T_141 ? 4'h2 : _T_2431; // @[Lookup.scala 33:37]
  wire [3:0] _T_2433 = _T_139 ? 4'h0 : _T_2432; // @[Lookup.scala 33:37]
  wire [3:0] _T_2434 = _T_137 ? 4'h0 : _T_2433; // @[Lookup.scala 33:37]
  wire [3:0] _T_2435 = _T_135 ? 4'h0 : _T_2434; // @[Lookup.scala 33:37]
  wire [3:0] _T_2436 = _T_133 ? 4'h7 : _T_2435; // @[Lookup.scala 33:37]
  wire [3:0] _T_2437 = _T_131 ? 4'h7 : _T_2436; // @[Lookup.scala 33:37]
  wire [3:0] rvcDestType = _T_129 ? 4'h7 : _T_2437; // @[Lookup.scala 33:37]
  wire  _T_2441 = 5'h4 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2443 = 5'h2 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2444 = 5'hf == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2445 = 5'h1 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2446 = 5'h6 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2447 = 5'h7 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2448 = 5'h0 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2450 = 5'h15 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2451 = 5'h17 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_2454 = 5'hc == instrType; // @[LookupTree.scala 24:34]
  wire  src1Type = _T_2446 | _T_2447 | _T_2448; // @[Mux.scala 27:72]
  wire  src2Type = _T_2441 | _T_2446 | _T_2447 | _T_2448 | _T_2450 | _T_2451 | _T_2454; // @[Mux.scala 27:72]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[IDU.scala 72:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[IDU.scala 72:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[IDU.scala 72:58]
  wire [4:0] rs2 = io_in_bits_instr[6:2]; // @[IDU.scala 75:24]
  wire  _T_2524 = 3'h0 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2525 = 3'h1 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2526 = 3'h2 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2527 = 3'h3 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2528 = 3'h4 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2529 = 3'h5 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2530 = 3'h6 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_2531 = 3'h7 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_2532 = _T_2524 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2533 = _T_2525 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2534 = _T_2526 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2535 = _T_2527 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2536 = _T_2528 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2537 = _T_2529 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2538 = _T_2530 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2539 = _T_2531 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2540 = _T_2532 | _T_2533; // @[Mux.scala 27:72]
  wire [3:0] _T_2541 = _T_2540 | _T_2534; // @[Mux.scala 27:72]
  wire [3:0] _T_2542 = _T_2541 | _T_2535; // @[Mux.scala 27:72]
  wire [3:0] _T_2543 = _T_2542 | _T_2536; // @[Mux.scala 27:72]
  wire [3:0] _T_2544 = _T_2543 | _T_2537; // @[Mux.scala 27:72]
  wire [3:0] _T_2545 = _T_2544 | _T_2538; // @[Mux.scala 27:72]
  wire [3:0] rs1p = _T_2545 | _T_2539; // @[Mux.scala 27:72]
  wire  _T_2548 = 3'h0 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2549 = 3'h1 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2550 = 3'h2 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2551 = 3'h3 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2552 = 3'h4 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2553 = 3'h5 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2554 = 3'h6 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_2555 = 3'h7 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_2556 = _T_2548 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2557 = _T_2549 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2558 = _T_2550 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2559 = _T_2551 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2560 = _T_2552 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2561 = _T_2553 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2562 = _T_2554 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2563 = _T_2555 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2564 = _T_2556 | _T_2557; // @[Mux.scala 27:72]
  wire [3:0] _T_2565 = _T_2564 | _T_2558; // @[Mux.scala 27:72]
  wire [3:0] _T_2566 = _T_2565 | _T_2559; // @[Mux.scala 27:72]
  wire [3:0] _T_2567 = _T_2566 | _T_2560; // @[Mux.scala 27:72]
  wire [3:0] _T_2568 = _T_2567 | _T_2561; // @[Mux.scala 27:72]
  wire [3:0] _T_2569 = _T_2568 | _T_2562; // @[Mux.scala 27:72]
  wire [3:0] rs2p = _T_2569 | _T_2563; // @[Mux.scala 27:72]
  wire [5:0] rvc_shamt = {io_in_bits_instr[12],rs2}; // @[Cat.scala 30:58]
  wire  _T_2574 = 4'h3 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2575 = 4'h1 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2576 = 4'h2 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2577 = 4'h4 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2578 = 4'h5 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2579 = 4'h6 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2580 = 4'h7 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2581 = 4'h8 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_2582 = 4'h9 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire [4:0] _T_2584 = _T_2574 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2585 = _T_2575 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2586 = _T_2576 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2587 = _T_2577 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2588 = _T_2578 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2589 = _T_2579 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2590 = _T_2580 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_2592 = _T_2582 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2594 = _T_2584 | _T_2585; // @[Mux.scala 27:72]
  wire [4:0] _T_2595 = _T_2594 | _T_2586; // @[Mux.scala 27:72]
  wire [4:0] _T_2596 = _T_2595 | _T_2587; // @[Mux.scala 27:72]
  wire [4:0] _T_2597 = _T_2596 | _T_2588; // @[Mux.scala 27:72]
  wire [4:0] _GEN_5 = {{1'd0}, _T_2589}; // @[Mux.scala 27:72]
  wire [4:0] _T_2598 = _T_2597 | _GEN_5; // @[Mux.scala 27:72]
  wire [4:0] _GEN_6 = {{1'd0}, _T_2590}; // @[Mux.scala 27:72]
  wire [4:0] _T_2599 = _T_2598 | _GEN_6; // @[Mux.scala 27:72]
  wire [4:0] _GEN_7 = {{4'd0}, _T_2581}; // @[Mux.scala 27:72]
  wire [4:0] _T_2600 = _T_2599 | _GEN_7; // @[Mux.scala 27:72]
  wire [4:0] _GEN_8 = {{3'd0}, _T_2592}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src1 = _T_2600 | _GEN_8; // @[Mux.scala 27:72]
  wire  _T_2603 = 3'h3 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_2604 = 3'h1 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_2605 = 3'h2 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_2606 = 3'h4 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_2607 = 3'h5 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_2608 = 3'h6 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_2609 = 3'h7 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire [3:0] _GEN_9 = {{1'd0}, rvcSrc2Type}; // @[LookupTree.scala 24:34]
  wire  _T_2610 = 4'h8 == _GEN_9; // @[LookupTree.scala 24:34]
  wire  _T_2611 = 4'h9 == _GEN_9; // @[LookupTree.scala 24:34]
  wire [4:0] _T_2613 = _T_2603 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2614 = _T_2604 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2615 = _T_2605 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2616 = _T_2606 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2617 = _T_2607 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2618 = _T_2608 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2619 = _T_2609 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_2621 = _T_2611 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2623 = _T_2613 | _T_2614; // @[Mux.scala 27:72]
  wire [4:0] _T_2624 = _T_2623 | _T_2615; // @[Mux.scala 27:72]
  wire [4:0] _T_2625 = _T_2624 | _T_2616; // @[Mux.scala 27:72]
  wire [4:0] _T_2626 = _T_2625 | _T_2617; // @[Mux.scala 27:72]
  wire [4:0] _GEN_11 = {{1'd0}, _T_2618}; // @[Mux.scala 27:72]
  wire [4:0] _T_2627 = _T_2626 | _GEN_11; // @[Mux.scala 27:72]
  wire [4:0] _GEN_12 = {{1'd0}, _T_2619}; // @[Mux.scala 27:72]
  wire [4:0] _T_2628 = _T_2627 | _GEN_12; // @[Mux.scala 27:72]
  wire [4:0] _GEN_13 = {{4'd0}, _T_2610}; // @[Mux.scala 27:72]
  wire [4:0] _T_2629 = _T_2628 | _GEN_13; // @[Mux.scala 27:72]
  wire [4:0] _GEN_14 = {{3'd0}, _T_2621}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src2 = _T_2629 | _GEN_14; // @[Mux.scala 27:72]
  wire  _T_2632 = 4'h3 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2633 = 4'h1 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2634 = 4'h2 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2635 = 4'h4 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2636 = 4'h5 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2637 = 4'h6 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2638 = 4'h7 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2639 = 4'h8 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_2640 = 4'h9 == rvcDestType; // @[LookupTree.scala 24:34]
  wire [4:0] _T_2642 = _T_2632 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2643 = _T_2633 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2644 = _T_2634 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2645 = _T_2635 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2646 = _T_2636 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2647 = _T_2637 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_2648 = _T_2638 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_2650 = _T_2640 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_2652 = _T_2642 | _T_2643; // @[Mux.scala 27:72]
  wire [4:0] _T_2653 = _T_2652 | _T_2644; // @[Mux.scala 27:72]
  wire [4:0] _T_2654 = _T_2653 | _T_2645; // @[Mux.scala 27:72]
  wire [4:0] _T_2655 = _T_2654 | _T_2646; // @[Mux.scala 27:72]
  wire [4:0] _GEN_15 = {{1'd0}, _T_2647}; // @[Mux.scala 27:72]
  wire [4:0] _T_2656 = _T_2655 | _GEN_15; // @[Mux.scala 27:72]
  wire [4:0] _GEN_16 = {{1'd0}, _T_2648}; // @[Mux.scala 27:72]
  wire [4:0] _T_2657 = _T_2656 | _GEN_16; // @[Mux.scala 27:72]
  wire [4:0] _GEN_17 = {{4'd0}, _T_2639}; // @[Mux.scala 27:72]
  wire [4:0] _T_2658 = _T_2657 | _GEN_17; // @[Mux.scala 27:72]
  wire [4:0] _GEN_18 = {{3'd0}, _T_2650}; // @[Mux.scala 27:72]
  wire [4:0] rvc_dest = _T_2658 | _GEN_18; // @[Mux.scala 27:72]
  wire  _T_2667 = io_in_bits_instr[14:12] == 3'h1 & io_in_bits_instr[6:0] == 7'h33 & io_in_bits_instr[26:25] == 2'h3; // @[IDU.scala 99:80]
  wire  src3fromhead = _T_2667 | io_in_bits_instr[26:25] == 2'h2 & io_in_bits_instr[14:12] == 3'h5 & io_in_bits_instr[6:
    0] == 7'h3b; // @[IDU.scala 100:21]
  wire  _T_2681 = io_in_bits_instr[14:12] == 3'h0; // @[IDU.scala 102:92]
  wire  insb = fuOpType == 7'h56 & io_in_bits_instr[24:23] == 2'h0 & io_in_bits_instr[14:12] == 3'h0; // @[IDU.scala 102:76]
  wire [4:0] rfSrc1 = isRVC ? rvc_src1 : rs; // @[IDU.scala 103:19]
  wire [4:0] rfSrc2 = isRVC ? rvc_src2 : rt; // @[IDU.scala 104:19]
  wire [4:0] rfDest = isRVC ? rvc_dest : rd; // @[IDU.scala 105:19]
  wire [4:0] _T_2692 = instrType == 5'h14 & fuOpType[6:1] == 6'h3f & _T_2681 | insb ? rd : 5'h0; // @[IDU.scala 106:79]
  wire [4:0] _T_2693 = instrType == 5'h1c ? rd : _T_2692; // @[IDU.scala 106:49]
  wire [51:0] _T_2704 = io_in_bits_instr[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2705 = {_T_2704,io_in_bits_instr[31:20]}; // @[Cat.scala 30:58]
  wire [11:0] _T_2708 = {io_in_bits_instr[31:25],rd}; // @[Cat.scala 30:58]
  wire [51:0] _T_2711 = _T_2708[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2712 = {_T_2711,io_in_bits_instr[31:25],rd}; // @[Cat.scala 30:58]
  wire [12:0] _T_2724 = {io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}; // @[Cat.scala 30:58]
  wire [50:0] _T_2727 = _T_2724[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2728 = {_T_2727,io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8]
    ,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_2730 = {io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_2733 = _T_2730[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2734 = {_T_2733,io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [20:0] _T_2739 = {io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0}
    ; // @[Cat.scala 30:58]
  wire [42:0] _T_2742 = _T_2739[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2743 = {_T_2742,io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:
    21],1'h0}; // @[Cat.scala 30:58]
  wire [57:0] _T_2747 = io_in_bits_instr[25] ? 58'h3ffffffffffffff : 58'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2748 = {_T_2747,io_in_bits_instr[25:20]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2755 = {47'h0,io_in_bits_instr[31:15]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2765 = _T_2441 ? _T_2705 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2766 = _T_2443 ? _T_2712 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2767 = _T_2444 ? _T_2712 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2768 = _T_2445 ? _T_2728 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2769 = _T_2446 ? _T_2734 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2770 = _T_2447 ? _T_2743 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2771 = _T_2450 ? _T_2748 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2772 = _T_2451 ? _T_2748 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2773 = _T_2454 ? _T_2755 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2774 = _T_2765 | _T_2766; // @[Mux.scala 27:72]
  wire [63:0] _T_2775 = _T_2774 | _T_2767; // @[Mux.scala 27:72]
  wire [63:0] _T_2776 = _T_2775 | _T_2768; // @[Mux.scala 27:72]
  wire [63:0] _T_2777 = _T_2776 | _T_2769; // @[Mux.scala 27:72]
  wire [63:0] _T_2778 = _T_2777 | _T_2770; // @[Mux.scala 27:72]
  wire [63:0] _T_2779 = _T_2778 | _T_2771; // @[Mux.scala 27:72]
  wire [63:0] _T_2780 = _T_2779 | _T_2772; // @[Mux.scala 27:72]
  wire [63:0] imm = _T_2780 | _T_2773; // @[Mux.scala 27:72]
  wire [63:0] _T_2786 = {56'h0,io_in_bits_instr[3:2],io_in_bits_instr[12],io_in_bits_instr[6:4],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_2791 = {55'h0,io_in_bits_instr[4:2],io_in_bits_instr[12],io_in_bits_instr[6:5],3'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_2795 = {56'h0,io_in_bits_instr[8:7],io_in_bits_instr[12:9],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_2799 = {55'h0,io_in_bits_instr[9:7],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_2804 = {57'h0,io_in_bits_instr[5],io_in_bits_instr[12:10],io_in_bits_instr[6],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_2808 = {56'h0,io_in_bits_instr[6:5],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 30:58]
  wire [11:0] _T_2826 = {io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],
    io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 30:58]
  wire [51:0] _T_2829 = _T_2826[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2830 = {_T_2829,io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],
    io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 30:58]
  wire [8:0] _T_2836 = {io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],
    io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 30:58]
  wire [54:0] _T_2839 = _T_2836[8] ? 55'h7fffffffffffff : 55'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2840 = {_T_2839,io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],
    io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 30:58]
  wire [57:0] _T_2846 = rvc_shamt[5] ? 58'h3ffffffffffffff : 58'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2847 = {_T_2846,io_in_bits_instr[12],rs2}; // @[Cat.scala 30:58]
  wire [17:0] _T_2850 = {io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 30:58]
  wire [45:0] _T_2853 = _T_2850[17] ? 46'h3fffffffffff : 46'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2854 = {_T_2853,io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 30:58]
  wire [9:0] _T_2867 = {io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],
    io_in_bits_instr[6],4'h0}; // @[Cat.scala 30:58]
  wire [53:0] _T_2870 = _T_2867[9] ? 54'h3fffffffffffff : 54'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2871 = {_T_2870,io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],
    io_in_bits_instr[6],4'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_2877 = {54'h0,io_in_bits_instr[10:7],io_in_bits_instr[12:11],io_in_bits_instr[5],io_in_bits_instr[6],2'h0
    }; // @[Cat.scala 30:58]
  wire  _T_2879 = 5'h0 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2880 = 5'h1 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2881 = 5'h2 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2882 = 5'h3 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2883 = 5'h4 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2884 = 5'h5 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2885 = 5'h6 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2886 = 5'h7 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2887 = 5'h8 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2888 = 5'h9 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2889 = 5'ha == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2890 = 5'hb == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2891 = 5'hc == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2892 = 5'hd == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2893 = 5'he == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_2894 = 5'hf == rvcImmType; // @[LookupTree.scala 24:34]
  wire [63:0] _T_2896 = _T_2879 ? _T_2786 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2897 = _T_2880 ? _T_2791 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2898 = _T_2881 ? _T_2795 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2899 = _T_2882 ? _T_2799 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2900 = _T_2883 ? _T_2804 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2901 = _T_2884 ? _T_2808 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2902 = _T_2885 ? _T_2804 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2903 = _T_2886 ? _T_2808 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2904 = _T_2887 ? _T_2830 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2905 = _T_2888 ? _T_2840 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2906 = _T_2889 ? _T_2847 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2907 = _T_2890 ? _T_2854 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2908 = _T_2891 ? _T_2847 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2909 = _T_2892 ? _T_2871 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2910 = _T_2893 ? _T_2877 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2911 = _T_2894 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_2913 = _T_2896 | _T_2897; // @[Mux.scala 27:72]
  wire [63:0] _T_2914 = _T_2913 | _T_2898; // @[Mux.scala 27:72]
  wire [63:0] _T_2915 = _T_2914 | _T_2899; // @[Mux.scala 27:72]
  wire [63:0] _T_2916 = _T_2915 | _T_2900; // @[Mux.scala 27:72]
  wire [63:0] _T_2917 = _T_2916 | _T_2901; // @[Mux.scala 27:72]
  wire [63:0] _T_2918 = _T_2917 | _T_2902; // @[Mux.scala 27:72]
  wire [63:0] _T_2919 = _T_2918 | _T_2903; // @[Mux.scala 27:72]
  wire [63:0] _T_2920 = _T_2919 | _T_2904; // @[Mux.scala 27:72]
  wire [63:0] _T_2921 = _T_2920 | _T_2905; // @[Mux.scala 27:72]
  wire [63:0] _T_2922 = _T_2921 | _T_2906; // @[Mux.scala 27:72]
  wire [63:0] _T_2923 = _T_2922 | _T_2907; // @[Mux.scala 27:72]
  wire [63:0] _T_2924 = _T_2923 | _T_2908; // @[Mux.scala 27:72]
  wire [63:0] _T_2925 = _T_2924 | _T_2909; // @[Mux.scala 27:72]
  wire [63:0] _T_2926 = _T_2925 | _T_2910; // @[Mux.scala 27:72]
  wire [63:0] immrvc = _T_2926 | _T_2911; // @[Mux.scala 27:72]
  wire  _T_2929 = fuType == 4'h0; // @[IDU.scala 151:16]
  wire  _T_2932 = rfDest == 5'h1 | rfDest == 5'h5; // @[IDU.scala 152:42]
  wire [6:0] _GEN_0 = _T_2932 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[IDU.scala 153:{57,85} 47:29]
  wire  _T_2938 = rfSrc1 == 5'h1 | rfSrc1 == 5'h5; // @[IDU.scala 152:42]
  wire [6:0] _GEN_1 = _T_2938 ? 7'h5e : _GEN_0; // @[IDU.scala 155:{29,57}]
  wire [6:0] _GEN_2 = _T_2932 ? 7'h5c : _GEN_1; // @[IDU.scala 156:{29,57}]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[IDU.scala 154:40]
  wire  _T_2956 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_2957 = ~hasIntr; // @[IDU.scala 181:51]
  wire [7:0] _T_3004 = {7'h17 == fuOpType,7'h16 == fuOpType,7'h15 == fuOpType,7'h14 == fuOpType,7'h11 == fuOpType,7'h10
     == fuOpType,7'h5a == fuOpType,7'h58 == fuOpType}; // @[IDU.scala 209:84]
  assign io_in_ready = ~io_in_valid | _T_2956 & ~hasIntr; // @[IDU.scala 181:31]
  assign io_out_valid = io_in_valid; // @[IDU.scala 180:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[IDU.scala 182:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[IDU.scala 182:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[IDU.scala 182:18]
  assign io_out_bits_cf_exceptionVec_1 = |io_in_bits_pc[38:32] & ~DTLBENABLE; // @[IDU.scala 200:98]
  assign io_out_bits_cf_exceptionVec_2 = instrType == 5'h0 & _T_2957 & io_in_valid; // @[IDU.scala 197:83]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[IDU.scala 198:47]
  assign io_out_bits_cf_intrVec_0 = intrVec[0]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_1 = intrVec[1]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_2 = intrVec[2]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_3 = intrVec[3]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_4 = intrVec[4]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_5 = intrVec[5]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_6 = intrVec[6]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_7 = intrVec[7]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_8 = intrVec[8]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_9 = intrVec[9]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_10 = intrVec[10]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_11 = intrVec[11]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[IDU.scala 182:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_bits_crossPageIPFFix; // @[IDU.scala 182:18]
  assign io_out_bits_cf_instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 5'h0 :
    decodeList_0; // @[IDU.scala 38:75]
  assign io_out_bits_ctrl_src1Type = io_in_bits_instr[6:0] == 7'h37 ? 1'h0 : src1Type; // @[IDU.scala 160:35]
  assign io_out_bits_ctrl_src2Type = _T_2441 | _T_2446 | _T_2447 | _T_2448 | _T_2450 | _T_2451 | _T_2454; // @[Mux.scala 27:72]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h1 :
    decodeList_1; // @[IDU.scala 38:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 4'h0 ? _GEN_3 : fuOpType; // @[IDU.scala 151:32 47:29]
  assign io_out_bits_ctrl_funct3 = io_in_bits_instr[14:12]; // @[IDU.scala 49:35]
  assign io_out_bits_ctrl_func24 = io_in_bits_instr[24]; // @[IDU.scala 50:35]
  assign io_out_bits_ctrl_func23 = io_in_bits_instr[23]; // @[IDU.scala 51:35]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rfSrc1; // @[IDU.scala 109:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rfSrc2 : 5'h0; // @[IDU.scala 110:33]
  assign io_out_bits_ctrl_rfSrc3 = src3fromhead ? io_in_bits_instr[31:27] : _T_2693; // @[IDU.scala 106:19]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[Decode.scala 39:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rfDest : 5'h0; // @[IDU.scala 113:33]
  assign io_out_bits_ctrl_isMou = fuType == 4'h8; // @[IDU.scala 206:36]
  assign io_out_bits_data_imm = isRVC ? immrvc : imm; // @[IDU.scala 149:31]
  assign io_isBranch = |_T_3004 & _T_2929; // @[IDU.scala 209:95]
endmodule
module Decoder_1(
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  input  [63:0] intrVecIDU
);
  wire [11:0] intrVec = intrVecIDU[11:0];
  assign io_out_bits_cf_intrVec_0 = intrVec[0]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_1 = intrVec[1]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_2 = intrVec[2]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_3 = intrVec[3]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_4 = intrVec[4]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_5 = intrVec[5]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_6 = intrVec[6]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_7 = intrVec[7]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_8 = intrVec[8]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_9 = intrVec[9]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_10 = intrVec[10]; // @[IDU.scala 190:38]
  assign io_out_bits_cf_intrVec_11 = intrVec[11]; // @[IDU.scala 190:38]
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_instr,
  input  [38:0] io_in_0_bits_pc,
  input  [38:0] io_in_0_bits_pnpc,
  input         io_in_0_bits_exceptionVec_12,
  input  [3:0]  io_in_0_bits_brIdx,
  input         io_in_0_bits_crossPageIPFFix,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [63:0] io_out_0_bits_cf_runahead_checkpoint_id,
  output [4:0]  io_out_0_bits_cf_instrType,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [3:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [2:0]  io_out_0_bits_ctrl_funct3,
  output        io_out_0_bits_ctrl_func24,
  output        io_out_0_bits_ctrl_func23,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output [4:0]  io_out_0_bits_ctrl_rfSrc3,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output        io_out_0_bits_ctrl_isMou,
  output [63:0] io_out_0_bits_data_imm,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  input         vmEnable,
  input  [63:0] intrVec
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  decoder1_io_in_ready; // @[IDU.scala 218:25]
  wire  decoder1_io_in_valid; // @[IDU.scala 218:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[IDU.scala 218:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[IDU.scala 218:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[IDU.scala 218:25]
  wire  decoder1_io_in_bits_exceptionVec_12; // @[IDU.scala 218:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[IDU.scala 218:25]
  wire  decoder1_io_in_bits_crossPageIPFFix; // @[IDU.scala 218:25]
  wire  decoder1_io_out_ready; // @[IDU.scala 218:25]
  wire  decoder1_io_out_valid; // @[IDU.scala 218:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[IDU.scala 218:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[IDU.scala 218:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 218:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 218:25]
  wire [4:0] decoder1_io_out_bits_cf_instrType; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 218:25]
  wire [3:0] decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 218:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 218:25]
  wire [2:0] decoder1_io_out_bits_ctrl_funct3; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_ctrl_func24; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_ctrl_func23; // @[IDU.scala 218:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 218:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 218:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc3; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 218:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 218:25]
  wire  decoder1_io_out_bits_ctrl_isMou; // @[IDU.scala 218:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[IDU.scala 218:25]
  wire  decoder1_io_isBranch; // @[IDU.scala 218:25]
  wire  decoder1_DTLBENABLE; // @[IDU.scala 218:25]
  wire [63:0] decoder1_intrVecIDU; // @[IDU.scala 218:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 219:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 219:25]
  wire [63:0] decoder2_intrVecIDU; // @[IDU.scala 219:25]
  wire  runahead_io_clock; // @[IDU.scala 233:24]
  wire [7:0] runahead_io_coreid; // @[IDU.scala 233:24]
  wire [7:0] runahead_io_index; // @[IDU.scala 233:24]
  wire  runahead_io_valid; // @[IDU.scala 233:24]
  wire  runahead_io_branch; // @[IDU.scala 233:24]
  wire  runahead_io_may_replay; // @[IDU.scala 233:24]
  wire [63:0] runahead_io_pc; // @[IDU.scala 233:24]
  wire [63:0] runahead_io_checkpoint_id; // @[IDU.scala 233:24]
  reg [63:0] checkpoint_id; // @[IDU.scala 230:30]
  wire [63:0] _T_3 = checkpoint_id + 64'h1; // @[IDU.scala 241:36]
  Decoder decoder1 ( // @[IDU.scala 218:25]
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder1_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder1_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder1_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder1_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_cf_instrType(decoder1_io_out_bits_cf_instrType),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_funct3(decoder1_io_out_bits_ctrl_funct3),
    .io_out_bits_ctrl_func24(decoder1_io_out_bits_ctrl_func24),
    .io_out_bits_ctrl_func23(decoder1_io_out_bits_ctrl_func23),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfSrc3(decoder1_io_out_bits_ctrl_rfSrc3),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isMou(decoder1_io_out_bits_ctrl_isMou),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .io_isBranch(decoder1_io_isBranch),
    .DTLBENABLE(decoder1_DTLBENABLE),
    .intrVecIDU(decoder1_intrVecIDU)
  );
  Decoder_1 decoder2 ( // @[IDU.scala 219:25]
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  DifftestRunaheadEvent runahead ( // @[IDU.scala 233:24]
    .io_clock(runahead_io_clock),
    .io_coreid(runahead_io_coreid),
    .io_index(runahead_io_index),
    .io_valid(runahead_io_valid),
    .io_branch(runahead_io_branch),
    .io_may_replay(runahead_io_may_replay),
    .io_pc(runahead_io_pc),
    .io_checkpoint_id(runahead_io_checkpoint_id)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[IDU.scala 220:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_crossPageIPFFix = decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 222:13]
  assign io_out_0_bits_cf_runahead_checkpoint_id = checkpoint_id; // @[IDU.scala 244:44]
  assign io_out_0_bits_cf_instrType = decoder1_io_out_bits_cf_instrType; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_funct3 = decoder1_io_out_bits_ctrl_funct3; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_func24 = decoder1_io_out_bits_ctrl_func24; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_func23 = decoder1_io_out_bits_ctrl_func23; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_rfSrc3 = decoder1_io_out_bits_ctrl_rfSrc3; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 222:13]
  assign io_out_0_bits_ctrl_isMou = decoder1_io_out_bits_ctrl_isMou; // @[IDU.scala 222:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[IDU.scala 222:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 223:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 223:13]
  assign decoder1_io_in_valid = io_in_0_valid; // @[IDU.scala 220:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[IDU.scala 220:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[IDU.scala 220:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[IDU.scala 220:12]
  assign decoder1_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[IDU.scala 220:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[IDU.scala 220:12]
  assign decoder1_io_in_bits_crossPageIPFFix = io_in_0_bits_crossPageIPFFix; // @[IDU.scala 220:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[IDU.scala 222:13]
  assign decoder1_DTLBENABLE = vmEnable;
  assign decoder1_intrVecIDU = intrVec;
  assign decoder2_intrVecIDU = intrVec;
  assign runahead_io_clock = clock; // @[IDU.scala 234:29]
  assign runahead_io_coreid = 8'h0; // @[IDU.scala 235:29]
  assign runahead_io_index = 8'h0;
  assign runahead_io_valid = io_out_0_ready & io_out_0_valid; // @[Decoupled.scala 40:37]
  assign runahead_io_branch = decoder1_io_isBranch; // @[IDU.scala 237:29]
  assign runahead_io_may_replay = 1'h0;
  assign runahead_io_pc = {{25'd0}, io_out_0_bits_cf_pc}; // @[IDU.scala 238:29]
  assign runahead_io_checkpoint_id = checkpoint_id; // @[IDU.scala 239:29]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 230:30]
      checkpoint_id <= 64'h0; // @[IDU.scala 230:30]
    end else if (runahead_io_valid & runahead_io_branch) begin // @[IDU.scala 240:49]
      checkpoint_id <= _T_3; // @[IDU.scala 241:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  checkpoint_id = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_instr,
  input  [38:0] io_enq_bits_pc,
  input  [38:0] io_enq_bits_pnpc,
  input         io_enq_bits_exceptionVec_12,
  input  [3:0]  io_enq_bits_brIdx,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_instr,
  output [38:0] io_deq_bits_pc,
  output [38:0] io_deq_bits_pnpc,
  output        io_deq_bits_exceptionVec_12,
  output [3:0]  io_deq_bits_brIdx,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] MEM_instr [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_instr_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_instr_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [63:0] MEM_instr_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [63:0] MEM_instr_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_instr_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_instr_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_instr_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [38:0] MEM_pc [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_pc_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pc_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pc_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pc_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pc_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_pc_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_pc_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [38:0] MEM_pnpc [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_pnpc_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pnpc_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pnpc_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pnpc_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pnpc_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_pnpc_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_pnpc_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg  MEM_exceptionVec_12 [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_exceptionVec_12_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_exceptionVec_12_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [3:0] MEM_brIdx [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_brIdx_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_brIdx_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [3:0] MEM_brIdx_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [3:0] MEM_brIdx_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_brIdx_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_brIdx_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_brIdx_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [1:0] value; // @[Counter.scala 60:40]
  reg [1:0] value_1; // @[Counter.scala 60:40]
  reg  REG; // @[FlushableQueue.scala 26:35]
  wire  _T = value == value_1; // @[FlushableQueue.scala 28:41]
  wire  _T_2 = _T & ~REG; // @[FlushableQueue.scala 29:33]
  wire  _T_3 = _T & REG; // @[FlushableQueue.scala 30:32]
  wire  _T_4 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _value_T_1 = value + 2'h1; // @[Counter.scala 76:24]
  wire [1:0] _value_T_3 = value_1 + 2'h1; // @[Counter.scala 76:24]
  assign MEM_instr_MPORT_1_en = 1'h1;
  assign MEM_instr_MPORT_1_addr = value_1;
  assign MEM_instr_MPORT_1_data = MEM_instr[MEM_instr_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_instr_MPORT_data = io_enq_bits_instr;
  assign MEM_instr_MPORT_addr = value;
  assign MEM_instr_MPORT_mask = 1'h1;
  assign MEM_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_pc_MPORT_1_en = 1'h1;
  assign MEM_pc_MPORT_1_addr = value_1;
  assign MEM_pc_MPORT_1_data = MEM_pc[MEM_pc_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_pc_MPORT_data = io_enq_bits_pc;
  assign MEM_pc_MPORT_addr = value;
  assign MEM_pc_MPORT_mask = 1'h1;
  assign MEM_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_pnpc_MPORT_1_en = 1'h1;
  assign MEM_pnpc_MPORT_1_addr = value_1;
  assign MEM_pnpc_MPORT_1_data = MEM_pnpc[MEM_pnpc_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_pnpc_MPORT_data = io_enq_bits_pnpc;
  assign MEM_pnpc_MPORT_addr = value;
  assign MEM_pnpc_MPORT_mask = 1'h1;
  assign MEM_pnpc_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_exceptionVec_12_MPORT_1_en = 1'h1;
  assign MEM_exceptionVec_12_MPORT_1_addr = value_1;
  assign MEM_exceptionVec_12_MPORT_1_data = MEM_exceptionVec_12[MEM_exceptionVec_12_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_exceptionVec_12_MPORT_data = io_enq_bits_exceptionVec_12;
  assign MEM_exceptionVec_12_MPORT_addr = value;
  assign MEM_exceptionVec_12_MPORT_mask = 1'h1;
  assign MEM_exceptionVec_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_brIdx_MPORT_1_en = 1'h1;
  assign MEM_brIdx_MPORT_1_addr = value_1;
  assign MEM_brIdx_MPORT_1_data = MEM_brIdx[MEM_brIdx_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_brIdx_MPORT_data = io_enq_bits_brIdx;
  assign MEM_brIdx_MPORT_addr = value;
  assign MEM_brIdx_MPORT_mask = 1'h1;
  assign MEM_brIdx_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_3; // @[FlushableQueue.scala 46:19]
  assign io_deq_valid = ~_T_2; // @[FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = MEM_instr_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_pc = MEM_pc_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_pnpc = MEM_pnpc_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_12 = MEM_exceptionVec_12_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_brIdx = MEM_brIdx_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  always @(posedge clock) begin
    if (MEM_instr_MPORT_en & MEM_instr_MPORT_mask) begin
      MEM_instr[MEM_instr_MPORT_addr] <= MEM_instr_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_pc_MPORT_en & MEM_pc_MPORT_mask) begin
      MEM_pc[MEM_pc_MPORT_addr] <= MEM_pc_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_pnpc_MPORT_en & MEM_pnpc_MPORT_mask) begin
      MEM_pnpc[MEM_pnpc_MPORT_addr] <= MEM_pnpc_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_exceptionVec_12_MPORT_en & MEM_exceptionVec_12_MPORT_mask) begin
      MEM_exceptionVec_12[MEM_exceptionVec_12_MPORT_addr] <= MEM_exceptionVec_12_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_brIdx_MPORT_en & MEM_brIdx_MPORT_mask) begin
      MEM_brIdx[MEM_brIdx_MPORT_addr] <= MEM_brIdx_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 2'h0; // @[Counter.scala 60:40]
    end else if (io_flush) begin // @[FlushableQueue.scala 62:19]
      value <= 2'h0; // @[FlushableQueue.scala 64:21]
    end else if (_T_4) begin // @[FlushableQueue.scala 34:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 2'h0; // @[Counter.scala 60:40]
    end else if (io_flush) begin // @[FlushableQueue.scala 62:19]
      value_1 <= 2'h0; // @[FlushableQueue.scala 65:21]
    end else if (_T_5) begin // @[FlushableQueue.scala 38:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[FlushableQueue.scala 26:35]
      REG <= 1'h0; // @[FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[FlushableQueue.scala 62:19]
      REG <= 1'h0; // @[FlushableQueue.scala 67:16]
    end else if (_T_4 != _T_5) begin // @[FlushableQueue.scala 41:28]
      REG <= _T_4; // @[FlushableQueue.scala 42:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_exceptionVec_12[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_brIdx[initvar] = _RAND_4[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  REG = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [86:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [86:0] io_imem_resp_bits_user,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [63:0] io_out_0_bits_cf_runahead_checkpoint_id,
  output [4:0]  io_out_0_bits_cf_instrType,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [3:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [2:0]  io_out_0_bits_ctrl_funct3,
  output        io_out_0_bits_ctrl_func24,
  output        io_out_0_bits_ctrl_func23,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output [4:0]  io_out_0_bits_ctrl_rfSrc3,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output        io_out_0_bits_ctrl_isMou,
  output [63:0] io_out_0_bits_data_imm,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  output [3:0]  io_flushVec,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  input         io_ipf,
  input         flushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         vmEnable,
  input  [63:0] intrVec,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[Frontend.scala 96:20]
  wire  ifu_reset; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_req_ready; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_req_valid; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Frontend.scala 96:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_resp_ready; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_resp_valid; // @[Frontend.scala 96:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Frontend.scala 96:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[Frontend.scala 96:20]
  wire  ifu_io_out_ready; // @[Frontend.scala 96:20]
  wire  ifu_io_out_valid; // @[Frontend.scala 96:20]
  wire [63:0] ifu_io_out_bits_instr; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_out_bits_pc; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[Frontend.scala 96:20]
  wire  ifu_io_out_bits_exceptionVec_12; // @[Frontend.scala 96:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_redirect_target; // @[Frontend.scala 96:20]
  wire  ifu_io_redirect_valid; // @[Frontend.scala 96:20]
  wire [3:0] ifu_io_flushVec; // @[Frontend.scala 96:20]
  wire  ifu_io_ipf; // @[Frontend.scala 96:20]
  wire  ifu_flushICache; // @[Frontend.scala 96:20]
  wire  ifu_bpuUpdateReq_valid; // @[Frontend.scala 96:20]
  wire [38:0] ifu_bpuUpdateReq_pc; // @[Frontend.scala 96:20]
  wire  ifu_bpuUpdateReq_isMissPredict; // @[Frontend.scala 96:20]
  wire [38:0] ifu_bpuUpdateReq_actualTarget; // @[Frontend.scala 96:20]
  wire  ifu_bpuUpdateReq_actualTaken; // @[Frontend.scala 96:20]
  wire [6:0] ifu_bpuUpdateReq_fuOpType; // @[Frontend.scala 96:20]
  wire [1:0] ifu_bpuUpdateReq_btbType; // @[Frontend.scala 96:20]
  wire  ifu_bpuUpdateReq_isRVC; // @[Frontend.scala 96:20]
  wire  ifu_flushTLB; // @[Frontend.scala 96:20]
  wire  ibf_clock; // @[Frontend.scala 97:19]
  wire  ibf_reset; // @[Frontend.scala 97:19]
  wire  ibf_io_in_ready; // @[Frontend.scala 97:19]
  wire  ibf_io_in_valid; // @[Frontend.scala 97:19]
  wire [63:0] ibf_io_in_bits_instr; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_in_bits_pc; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[Frontend.scala 97:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[Frontend.scala 97:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[Frontend.scala 97:19]
  wire  ibf_io_out_ready; // @[Frontend.scala 97:19]
  wire  ibf_io_out_valid; // @[Frontend.scala 97:19]
  wire [63:0] ibf_io_out_bits_instr; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_out_bits_pc; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[Frontend.scala 97:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[Frontend.scala 97:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[Frontend.scala 97:19]
  wire  ibf_io_out_bits_crossPageIPFFix; // @[Frontend.scala 97:19]
  wire  ibf_io_flush; // @[Frontend.scala 97:19]
  wire  idu_clock; // @[Frontend.scala 98:20]
  wire  idu_reset; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_ready; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_valid; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_bits_crossPageIPFFix; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_ready; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_valid; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_cf_instrType; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 98:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 98:20]
  wire [2:0] idu_io_out_0_bits_ctrl_funct3; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_func24; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_func23; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc3; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_isMou; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 98:20]
  wire  idu_vmEnable; // @[Frontend.scala 98:20]
  wire [63:0] idu_intrVec; // @[Frontend.scala 98:20]
  wire  FlushableQueue_clock; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_reset; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_enq_valid; // @[FlushableQueue.scala 94:21]
  wire [63:0] FlushableQueue_io_enq_bits_instr; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_enq_bits_pc; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_enq_bits_pnpc; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 94:21]
  wire [3:0] FlushableQueue_io_enq_bits_brIdx; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_deq_ready; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_deq_valid; // @[FlushableQueue.scala 94:21]
  wire [63:0] FlushableQueue_io_deq_bits_instr; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_deq_bits_pc; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_deq_bits_pnpc; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_deq_bits_exceptionVec_12; // @[FlushableQueue.scala 94:21]
  wire [3:0] FlushableQueue_io_deq_bits_brIdx; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_flush; // @[FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [63:0] r_instr; // @[Reg.scala 15:16]
  reg [38:0] r_pc; // @[Reg.scala 15:16]
  reg [38:0] r_pnpc; // @[Reg.scala 15:16]
  reg  r_exceptionVec_12; // @[Reg.scala 15:16]
  reg [3:0] r_brIdx; // @[Reg.scala 15:16]
  reg  r_crossPageIPFFix; // @[Reg.scala 15:16]
  IFU_inorder ifu ( // @[Frontend.scala 96:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ifu_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_ipf(ifu_io_ipf),
    .flushICache(ifu_flushICache),
    .bpuUpdateReq_valid(ifu_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(ifu_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(ifu_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(ifu_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(ifu_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(ifu_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(ifu_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(ifu_bpuUpdateReq_isRVC),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[Frontend.scala 97:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossPageIPFFix(ibf_io_out_bits_crossPageIPFFix),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[Frontend.scala 98:20]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossPageIPFFix(idu_io_in_0_bits_crossPageIPFFix),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(idu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_runahead_checkpoint_id(idu_io_out_0_bits_cf_runahead_checkpoint_id),
    .io_out_0_bits_cf_instrType(idu_io_out_0_bits_cf_instrType),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_funct3(idu_io_out_0_bits_ctrl_funct3),
    .io_out_0_bits_ctrl_func24(idu_io_out_0_bits_ctrl_func24),
    .io_out_0_bits_ctrl_func23(idu_io_out_0_bits_ctrl_func23),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfSrc3(idu_io_out_0_bits_ctrl_rfSrc3),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isMou(idu_io_out_0_bits_ctrl_isMou),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    .vmEnable(idu_vmEnable),
    .intrVec(idu_intrVec)
  );
  FlushableQueue FlushableQueue ( // @[FlushableQueue.scala 94:21]
    .clock(FlushableQueue_clock),
    .reset(FlushableQueue_reset),
    .io_enq_ready(FlushableQueue_io_enq_ready),
    .io_enq_valid(FlushableQueue_io_enq_valid),
    .io_enq_bits_instr(FlushableQueue_io_enq_bits_instr),
    .io_enq_bits_pc(FlushableQueue_io_enq_bits_pc),
    .io_enq_bits_pnpc(FlushableQueue_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_12(FlushableQueue_io_enq_bits_exceptionVec_12),
    .io_enq_bits_brIdx(FlushableQueue_io_enq_bits_brIdx),
    .io_deq_ready(FlushableQueue_io_deq_ready),
    .io_deq_valid(FlushableQueue_io_deq_valid),
    .io_deq_bits_instr(FlushableQueue_io_deq_bits_instr),
    .io_deq_bits_pc(FlushableQueue_io_deq_bits_pc),
    .io_deq_bits_pnpc(FlushableQueue_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_12(FlushableQueue_io_deq_bits_exceptionVec_12),
    .io_deq_bits_brIdx(FlushableQueue_io_deq_bits_brIdx),
    .io_flush(FlushableQueue_io_flush)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[Frontend.scala 118:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Frontend.scala 118:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[Frontend.scala 118:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[Frontend.scala 118:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_crossPageIPFFix = idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_runahead_checkpoint_id = idu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Frontend.scala 113:10]
  assign io_out_0_bits_cf_instrType = idu_io_out_0_bits_cf_instrType; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_funct3 = idu_io_out_0_bits_ctrl_funct3; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_func24 = idu_io_out_0_bits_ctrl_func24; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_func23 = idu_io_out_0_bits_ctrl_func23; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_rfSrc3 = idu_io_out_0_bits_ctrl_rfSrc3; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 113:10]
  assign io_out_0_bits_ctrl_isMou = idu_io_out_0_bits_ctrl_isMou; // @[Frontend.scala 113:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 113:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 113:10]
  assign io_flushVec = ifu_io_flushVec; // @[Frontend.scala 115:15]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[Frontend.scala 118:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[Frontend.scala 118:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Frontend.scala 118:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[Frontend.scala 118:11]
  assign ifu_io_out_ready = FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[Frontend.scala 114:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[Frontend.scala 114:15]
  assign ifu_io_ipf = io_ipf; // @[Frontend.scala 117:10]
  assign ifu_flushICache = flushICache;
  assign ifu_bpuUpdateReq_valid = bpuUpdateReq_valid;
  assign ifu_bpuUpdateReq_pc = bpuUpdateReq_pc;
  assign ifu_bpuUpdateReq_isMissPredict = bpuUpdateReq_isMissPredict;
  assign ifu_bpuUpdateReq_actualTarget = bpuUpdateReq_actualTarget;
  assign ifu_bpuUpdateReq_actualTaken = bpuUpdateReq_actualTaken;
  assign ifu_bpuUpdateReq_fuOpType = bpuUpdateReq_fuOpType;
  assign ifu_bpuUpdateReq_btbType = bpuUpdateReq_btbType;
  assign ifu_bpuUpdateReq_isRVC = bpuUpdateReq_isRVC;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = FlushableQueue_io_deq_valid; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_instr = FlushableQueue_io_deq_bits_instr; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_pc = FlushableQueue_io_deq_bits_pc; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_pnpc = FlushableQueue_io_deq_bits_pnpc; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_exceptionVec_12 = FlushableQueue_io_deq_bits_exceptionVec_12; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_brIdx = FlushableQueue_io_deq_bits_brIdx; // @[Frontend.scala 104:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[Frontend.scala 112:34]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_0_valid = REG; // @[Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = r_instr; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = r_pc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = r_pnpc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = r_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = r_brIdx; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossPageIPFFix = r_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[Frontend.scala 113:10]
  assign idu_vmEnable = vmEnable;
  assign idu_intrVec = intrVec;
  assign FlushableQueue_clock = clock;
  assign FlushableQueue_reset = reset;
  assign FlushableQueue_io_enq_valid = ifu_io_out_valid; // @[FlushableQueue.scala 95:22]
  assign FlushableQueue_io_enq_bits_instr = ifu_io_out_bits_instr; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_pc = ifu_io_out_bits_pc; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_exceptionVec_12 = ifu_io_out_bits_exceptionVec_12; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_deq_ready = ibf_io_in_ready; // @[Frontend.scala 104:11]
  assign FlushableQueue_io_flush = ifu_io_flushVec[0]; // @[Frontend.scala 107:58]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_instr <= ibf_io_out_bits_instr; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_pc <= ibf_io_out_bits_pc; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_pnpc <= ibf_io_out_bits_pnpc; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_brIdx <= ibf_io_out_bits_brIdx; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_crossPageIPFFix <= ibf_io_out_bits_crossPageIPFFix; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  r_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  r_exceptionVec_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_brIdx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  r_crossPageIPFFix = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstBoard(
  input        clock,
  input        reset,
  input        io_Wen_1,
  input        io_Wen_2,
  input        io_Wen_3,
  input        io_Wen_4,
  input        io_Wen_5,
  input        io_Wen_6,
  input        io_Wen_7,
  input        io_Wen_8,
  input        io_Wen_9,
  input        io_Wen_10,
  input        io_Wen_11,
  input        io_Wen_12,
  input        io_Wen_13,
  input        io_Wen_14,
  input        io_Wen_15,
  input        io_Wen_16,
  input        io_Wen_17,
  input        io_Wen_18,
  input        io_Wen_19,
  input        io_Wen_20,
  input        io_Wen_21,
  input        io_Wen_22,
  input        io_Wen_23,
  input        io_Wen_24,
  input        io_Wen_25,
  input        io_Wen_26,
  input        io_Wen_27,
  input        io_Wen_28,
  input        io_Wen_29,
  input        io_Wen_30,
  input        io_Wen_31,
  input        io_clear_1,
  input        io_clear_2,
  input        io_clear_3,
  input        io_clear_4,
  input        io_clear_5,
  input        io_clear_6,
  input        io_clear_7,
  input        io_clear_8,
  input        io_clear_9,
  input        io_clear_10,
  input        io_clear_11,
  input        io_clear_12,
  input        io_clear_13,
  input        io_clear_14,
  input        io_clear_15,
  input        io_clear_16,
  input        io_clear_17,
  input        io_clear_18,
  input        io_clear_19,
  input        io_clear_20,
  input        io_clear_21,
  input        io_clear_22,
  input        io_clear_23,
  input        io_clear_24,
  input        io_clear_25,
  input        io_clear_26,
  input        io_clear_27,
  input        io_clear_28,
  input        io_clear_29,
  input        io_clear_30,
  input        io_clear_31,
  input  [4:0] io_WInstNo_1,
  input  [4:0] io_WInstNo_2,
  input  [4:0] io_WInstNo_3,
  input  [4:0] io_WInstNo_4,
  input  [4:0] io_WInstNo_5,
  input  [4:0] io_WInstNo_6,
  input  [4:0] io_WInstNo_7,
  input  [4:0] io_WInstNo_8,
  input  [4:0] io_WInstNo_9,
  input  [4:0] io_WInstNo_10,
  input  [4:0] io_WInstNo_11,
  input  [4:0] io_WInstNo_12,
  input  [4:0] io_WInstNo_13,
  input  [4:0] io_WInstNo_14,
  input  [4:0] io_WInstNo_15,
  input  [4:0] io_WInstNo_16,
  input  [4:0] io_WInstNo_17,
  input  [4:0] io_WInstNo_18,
  input  [4:0] io_WInstNo_19,
  input  [4:0] io_WInstNo_20,
  input  [4:0] io_WInstNo_21,
  input  [4:0] io_WInstNo_22,
  input  [4:0] io_WInstNo_23,
  input  [4:0] io_WInstNo_24,
  input  [4:0] io_WInstNo_25,
  input  [4:0] io_WInstNo_26,
  input  [4:0] io_WInstNo_27,
  input  [4:0] io_WInstNo_28,
  input  [4:0] io_WInstNo_29,
  input  [4:0] io_WInstNo_30,
  input  [4:0] io_WInstNo_31,
  output       io_valid_1,
  output       io_valid_2,
  output       io_valid_3,
  output       io_valid_4,
  output       io_valid_5,
  output       io_valid_6,
  output       io_valid_7,
  output       io_valid_8,
  output       io_valid_9,
  output       io_valid_10,
  output       io_valid_11,
  output       io_valid_12,
  output       io_valid_13,
  output       io_valid_14,
  output       io_valid_15,
  output       io_valid_16,
  output       io_valid_17,
  output       io_valid_18,
  output       io_valid_19,
  output       io_valid_20,
  output       io_valid_21,
  output       io_valid_22,
  output       io_valid_23,
  output       io_valid_24,
  output       io_valid_25,
  output       io_valid_26,
  output       io_valid_27,
  output       io_valid_28,
  output       io_valid_29,
  output       io_valid_30,
  output       io_valid_31,
  output [4:0] io_RInstNo_1,
  output [4:0] io_RInstNo_2,
  output [4:0] io_RInstNo_3,
  output [4:0] io_RInstNo_4,
  output [4:0] io_RInstNo_5,
  output [4:0] io_RInstNo_6,
  output [4:0] io_RInstNo_7,
  output [4:0] io_RInstNo_8,
  output [4:0] io_RInstNo_9,
  output [4:0] io_RInstNo_10,
  output [4:0] io_RInstNo_11,
  output [4:0] io_RInstNo_12,
  output [4:0] io_RInstNo_13,
  output [4:0] io_RInstNo_14,
  output [4:0] io_RInstNo_15,
  output [4:0] io_RInstNo_16,
  output [4:0] io_RInstNo_17,
  output [4:0] io_RInstNo_18,
  output [4:0] io_RInstNo_19,
  output [4:0] io_RInstNo_20,
  output [4:0] io_RInstNo_21,
  output [4:0] io_RInstNo_22,
  output [4:0] io_RInstNo_23,
  output [4:0] io_RInstNo_24,
  output [4:0] io_RInstNo_25,
  output [4:0] io_RInstNo_26,
  output [4:0] io_RInstNo_27,
  output [4:0] io_RInstNo_28,
  output [4:0] io_RInstNo_29,
  output [4:0] io_RInstNo_30,
  output [4:0] io_RInstNo_31,
  input        io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
`endif // RANDOMIZE_REG_INIT
  reg  validBoard_1; // @[RF.scala 134:23]
  reg  validBoard_2; // @[RF.scala 134:23]
  reg  validBoard_3; // @[RF.scala 134:23]
  reg  validBoard_4; // @[RF.scala 134:23]
  reg  validBoard_5; // @[RF.scala 134:23]
  reg  validBoard_6; // @[RF.scala 134:23]
  reg  validBoard_7; // @[RF.scala 134:23]
  reg  validBoard_8; // @[RF.scala 134:23]
  reg  validBoard_9; // @[RF.scala 134:23]
  reg  validBoard_10; // @[RF.scala 134:23]
  reg  validBoard_11; // @[RF.scala 134:23]
  reg  validBoard_12; // @[RF.scala 134:23]
  reg  validBoard_13; // @[RF.scala 134:23]
  reg  validBoard_14; // @[RF.scala 134:23]
  reg  validBoard_15; // @[RF.scala 134:23]
  reg  validBoard_16; // @[RF.scala 134:23]
  reg  validBoard_17; // @[RF.scala 134:23]
  reg  validBoard_18; // @[RF.scala 134:23]
  reg  validBoard_19; // @[RF.scala 134:23]
  reg  validBoard_20; // @[RF.scala 134:23]
  reg  validBoard_21; // @[RF.scala 134:23]
  reg  validBoard_22; // @[RF.scala 134:23]
  reg  validBoard_23; // @[RF.scala 134:23]
  reg  validBoard_24; // @[RF.scala 134:23]
  reg  validBoard_25; // @[RF.scala 134:23]
  reg  validBoard_26; // @[RF.scala 134:23]
  reg  validBoard_27; // @[RF.scala 134:23]
  reg  validBoard_28; // @[RF.scala 134:23]
  reg  validBoard_29; // @[RF.scala 134:23]
  reg  validBoard_30; // @[RF.scala 134:23]
  reg  validBoard_31; // @[RF.scala 134:23]
  reg [4:0] InstBoard_1; // @[RF.scala 135:23]
  reg [4:0] InstBoard_2; // @[RF.scala 135:23]
  reg [4:0] InstBoard_3; // @[RF.scala 135:23]
  reg [4:0] InstBoard_4; // @[RF.scala 135:23]
  reg [4:0] InstBoard_5; // @[RF.scala 135:23]
  reg [4:0] InstBoard_6; // @[RF.scala 135:23]
  reg [4:0] InstBoard_7; // @[RF.scala 135:23]
  reg [4:0] InstBoard_8; // @[RF.scala 135:23]
  reg [4:0] InstBoard_9; // @[RF.scala 135:23]
  reg [4:0] InstBoard_10; // @[RF.scala 135:23]
  reg [4:0] InstBoard_11; // @[RF.scala 135:23]
  reg [4:0] InstBoard_12; // @[RF.scala 135:23]
  reg [4:0] InstBoard_13; // @[RF.scala 135:23]
  reg [4:0] InstBoard_14; // @[RF.scala 135:23]
  reg [4:0] InstBoard_15; // @[RF.scala 135:23]
  reg [4:0] InstBoard_16; // @[RF.scala 135:23]
  reg [4:0] InstBoard_17; // @[RF.scala 135:23]
  reg [4:0] InstBoard_18; // @[RF.scala 135:23]
  reg [4:0] InstBoard_19; // @[RF.scala 135:23]
  reg [4:0] InstBoard_20; // @[RF.scala 135:23]
  reg [4:0] InstBoard_21; // @[RF.scala 135:23]
  reg [4:0] InstBoard_22; // @[RF.scala 135:23]
  reg [4:0] InstBoard_23; // @[RF.scala 135:23]
  reg [4:0] InstBoard_24; // @[RF.scala 135:23]
  reg [4:0] InstBoard_25; // @[RF.scala 135:23]
  reg [4:0] InstBoard_26; // @[RF.scala 135:23]
  reg [4:0] InstBoard_27; // @[RF.scala 135:23]
  reg [4:0] InstBoard_28; // @[RF.scala 135:23]
  reg [4:0] InstBoard_29; // @[RF.scala 135:23]
  reg [4:0] InstBoard_30; // @[RF.scala 135:23]
  reg [4:0] InstBoard_31; // @[RF.scala 135:23]
  wire  _GEN_0 = io_clear_1 ? 1'h0 : validBoard_1; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_2 = io_Wen_1 | _GEN_0; // @[RF.scala 144:22 146:22]
  wire  _GEN_3 = io_clear_2 ? 1'h0 : validBoard_2; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_5 = io_Wen_2 | _GEN_3; // @[RF.scala 144:22 146:22]
  wire  _GEN_6 = io_clear_3 ? 1'h0 : validBoard_3; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_8 = io_Wen_3 | _GEN_6; // @[RF.scala 144:22 146:22]
  wire  _GEN_9 = io_clear_4 ? 1'h0 : validBoard_4; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_11 = io_Wen_4 | _GEN_9; // @[RF.scala 144:22 146:22]
  wire  _GEN_12 = io_clear_5 ? 1'h0 : validBoard_5; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_14 = io_Wen_5 | _GEN_12; // @[RF.scala 144:22 146:22]
  wire  _GEN_15 = io_clear_6 ? 1'h0 : validBoard_6; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_17 = io_Wen_6 | _GEN_15; // @[RF.scala 144:22 146:22]
  wire  _GEN_18 = io_clear_7 ? 1'h0 : validBoard_7; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_20 = io_Wen_7 | _GEN_18; // @[RF.scala 144:22 146:22]
  wire  _GEN_21 = io_clear_8 ? 1'h0 : validBoard_8; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_23 = io_Wen_8 | _GEN_21; // @[RF.scala 144:22 146:22]
  wire  _GEN_24 = io_clear_9 ? 1'h0 : validBoard_9; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_26 = io_Wen_9 | _GEN_24; // @[RF.scala 144:22 146:22]
  wire  _GEN_27 = io_clear_10 ? 1'h0 : validBoard_10; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_29 = io_Wen_10 | _GEN_27; // @[RF.scala 144:22 146:22]
  wire  _GEN_30 = io_clear_11 ? 1'h0 : validBoard_11; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_32 = io_Wen_11 | _GEN_30; // @[RF.scala 144:22 146:22]
  wire  _GEN_33 = io_clear_12 ? 1'h0 : validBoard_12; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_35 = io_Wen_12 | _GEN_33; // @[RF.scala 144:22 146:22]
  wire  _GEN_36 = io_clear_13 ? 1'h0 : validBoard_13; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_38 = io_Wen_13 | _GEN_36; // @[RF.scala 144:22 146:22]
  wire  _GEN_39 = io_clear_14 ? 1'h0 : validBoard_14; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_41 = io_Wen_14 | _GEN_39; // @[RF.scala 144:22 146:22]
  wire  _GEN_42 = io_clear_15 ? 1'h0 : validBoard_15; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_44 = io_Wen_15 | _GEN_42; // @[RF.scala 144:22 146:22]
  wire  _GEN_45 = io_clear_16 ? 1'h0 : validBoard_16; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_47 = io_Wen_16 | _GEN_45; // @[RF.scala 144:22 146:22]
  wire  _GEN_48 = io_clear_17 ? 1'h0 : validBoard_17; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_50 = io_Wen_17 | _GEN_48; // @[RF.scala 144:22 146:22]
  wire  _GEN_51 = io_clear_18 ? 1'h0 : validBoard_18; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_53 = io_Wen_18 | _GEN_51; // @[RF.scala 144:22 146:22]
  wire  _GEN_54 = io_clear_19 ? 1'h0 : validBoard_19; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_56 = io_Wen_19 | _GEN_54; // @[RF.scala 144:22 146:22]
  wire  _GEN_57 = io_clear_20 ? 1'h0 : validBoard_20; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_59 = io_Wen_20 | _GEN_57; // @[RF.scala 144:22 146:22]
  wire  _GEN_60 = io_clear_21 ? 1'h0 : validBoard_21; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_62 = io_Wen_21 | _GEN_60; // @[RF.scala 144:22 146:22]
  wire  _GEN_63 = io_clear_22 ? 1'h0 : validBoard_22; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_65 = io_Wen_22 | _GEN_63; // @[RF.scala 144:22 146:22]
  wire  _GEN_66 = io_clear_23 ? 1'h0 : validBoard_23; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_68 = io_Wen_23 | _GEN_66; // @[RF.scala 144:22 146:22]
  wire  _GEN_69 = io_clear_24 ? 1'h0 : validBoard_24; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_71 = io_Wen_24 | _GEN_69; // @[RF.scala 144:22 146:22]
  wire  _GEN_72 = io_clear_25 ? 1'h0 : validBoard_25; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_74 = io_Wen_25 | _GEN_72; // @[RF.scala 144:22 146:22]
  wire  _GEN_75 = io_clear_26 ? 1'h0 : validBoard_26; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_77 = io_Wen_26 | _GEN_75; // @[RF.scala 144:22 146:22]
  wire  _GEN_78 = io_clear_27 ? 1'h0 : validBoard_27; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_80 = io_Wen_27 | _GEN_78; // @[RF.scala 144:22 146:22]
  wire  _GEN_81 = io_clear_28 ? 1'h0 : validBoard_28; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_83 = io_Wen_28 | _GEN_81; // @[RF.scala 144:22 146:22]
  wire  _GEN_84 = io_clear_29 ? 1'h0 : validBoard_29; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_86 = io_Wen_29 | _GEN_84; // @[RF.scala 144:22 146:22]
  wire  _GEN_87 = io_clear_30 ? 1'h0 : validBoard_30; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_89 = io_Wen_30 | _GEN_87; // @[RF.scala 144:22 146:22]
  wire  _GEN_90 = io_clear_31 ? 1'h0 : validBoard_31; // @[RF.scala 134:23 147:30 148:23]
  wire  _GEN_92 = io_Wen_31 | _GEN_90; // @[RF.scala 144:22 146:22]
  assign io_valid_1 = validBoard_1; // @[RF.scala 159:13]
  assign io_valid_2 = validBoard_2; // @[RF.scala 159:13]
  assign io_valid_3 = validBoard_3; // @[RF.scala 159:13]
  assign io_valid_4 = validBoard_4; // @[RF.scala 159:13]
  assign io_valid_5 = validBoard_5; // @[RF.scala 159:13]
  assign io_valid_6 = validBoard_6; // @[RF.scala 159:13]
  assign io_valid_7 = validBoard_7; // @[RF.scala 159:13]
  assign io_valid_8 = validBoard_8; // @[RF.scala 159:13]
  assign io_valid_9 = validBoard_9; // @[RF.scala 159:13]
  assign io_valid_10 = validBoard_10; // @[RF.scala 159:13]
  assign io_valid_11 = validBoard_11; // @[RF.scala 159:13]
  assign io_valid_12 = validBoard_12; // @[RF.scala 159:13]
  assign io_valid_13 = validBoard_13; // @[RF.scala 159:13]
  assign io_valid_14 = validBoard_14; // @[RF.scala 159:13]
  assign io_valid_15 = validBoard_15; // @[RF.scala 159:13]
  assign io_valid_16 = validBoard_16; // @[RF.scala 159:13]
  assign io_valid_17 = validBoard_17; // @[RF.scala 159:13]
  assign io_valid_18 = validBoard_18; // @[RF.scala 159:13]
  assign io_valid_19 = validBoard_19; // @[RF.scala 159:13]
  assign io_valid_20 = validBoard_20; // @[RF.scala 159:13]
  assign io_valid_21 = validBoard_21; // @[RF.scala 159:13]
  assign io_valid_22 = validBoard_22; // @[RF.scala 159:13]
  assign io_valid_23 = validBoard_23; // @[RF.scala 159:13]
  assign io_valid_24 = validBoard_24; // @[RF.scala 159:13]
  assign io_valid_25 = validBoard_25; // @[RF.scala 159:13]
  assign io_valid_26 = validBoard_26; // @[RF.scala 159:13]
  assign io_valid_27 = validBoard_27; // @[RF.scala 159:13]
  assign io_valid_28 = validBoard_28; // @[RF.scala 159:13]
  assign io_valid_29 = validBoard_29; // @[RF.scala 159:13]
  assign io_valid_30 = validBoard_30; // @[RF.scala 159:13]
  assign io_valid_31 = validBoard_31; // @[RF.scala 159:13]
  assign io_RInstNo_1 = InstBoard_1; // @[RF.scala 160:13]
  assign io_RInstNo_2 = InstBoard_2; // @[RF.scala 160:13]
  assign io_RInstNo_3 = InstBoard_3; // @[RF.scala 160:13]
  assign io_RInstNo_4 = InstBoard_4; // @[RF.scala 160:13]
  assign io_RInstNo_5 = InstBoard_5; // @[RF.scala 160:13]
  assign io_RInstNo_6 = InstBoard_6; // @[RF.scala 160:13]
  assign io_RInstNo_7 = InstBoard_7; // @[RF.scala 160:13]
  assign io_RInstNo_8 = InstBoard_8; // @[RF.scala 160:13]
  assign io_RInstNo_9 = InstBoard_9; // @[RF.scala 160:13]
  assign io_RInstNo_10 = InstBoard_10; // @[RF.scala 160:13]
  assign io_RInstNo_11 = InstBoard_11; // @[RF.scala 160:13]
  assign io_RInstNo_12 = InstBoard_12; // @[RF.scala 160:13]
  assign io_RInstNo_13 = InstBoard_13; // @[RF.scala 160:13]
  assign io_RInstNo_14 = InstBoard_14; // @[RF.scala 160:13]
  assign io_RInstNo_15 = InstBoard_15; // @[RF.scala 160:13]
  assign io_RInstNo_16 = InstBoard_16; // @[RF.scala 160:13]
  assign io_RInstNo_17 = InstBoard_17; // @[RF.scala 160:13]
  assign io_RInstNo_18 = InstBoard_18; // @[RF.scala 160:13]
  assign io_RInstNo_19 = InstBoard_19; // @[RF.scala 160:13]
  assign io_RInstNo_20 = InstBoard_20; // @[RF.scala 160:13]
  assign io_RInstNo_21 = InstBoard_21; // @[RF.scala 160:13]
  assign io_RInstNo_22 = InstBoard_22; // @[RF.scala 160:13]
  assign io_RInstNo_23 = InstBoard_23; // @[RF.scala 160:13]
  assign io_RInstNo_24 = InstBoard_24; // @[RF.scala 160:13]
  assign io_RInstNo_25 = InstBoard_25; // @[RF.scala 160:13]
  assign io_RInstNo_26 = InstBoard_26; // @[RF.scala 160:13]
  assign io_RInstNo_27 = InstBoard_27; // @[RF.scala 160:13]
  assign io_RInstNo_28 = InstBoard_28; // @[RF.scala 160:13]
  assign io_RInstNo_29 = InstBoard_29; // @[RF.scala 160:13]
  assign io_RInstNo_30 = InstBoard_30; // @[RF.scala 160:13]
  assign io_RInstNo_31 = InstBoard_31; // @[RF.scala 160:13]
  always @(posedge clock) begin
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_1 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_1 <= _GEN_2;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_2 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_2 <= _GEN_5;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_3 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_3 <= _GEN_8;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_4 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_4 <= _GEN_11;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_5 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_5 <= _GEN_14;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_6 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_6 <= _GEN_17;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_7 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_7 <= _GEN_20;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_8 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_8 <= _GEN_23;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_9 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_9 <= _GEN_26;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_10 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_10 <= _GEN_29;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_11 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_11 <= _GEN_32;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_12 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_12 <= _GEN_35;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_13 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_13 <= _GEN_38;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_14 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_14 <= _GEN_41;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_15 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_15 <= _GEN_44;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_16 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_16 <= _GEN_47;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_17 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_17 <= _GEN_50;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_18 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_18 <= _GEN_53;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_19 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_19 <= _GEN_56;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_20 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_20 <= _GEN_59;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_21 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_21 <= _GEN_62;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_22 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_22 <= _GEN_65;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_23 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_23 <= _GEN_68;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_24 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_24 <= _GEN_71;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_25 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_25 <= _GEN_74;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_26 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_26 <= _GEN_77;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_27 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_27 <= _GEN_80;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_28 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_28 <= _GEN_83;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_29 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_29 <= _GEN_86;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_30 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_30 <= _GEN_89;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      validBoard_31 <= 1'h0; // @[RF.scala 138:21]
    end else begin
      validBoard_31 <= _GEN_92;
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_1 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_1) begin // @[RF.scala 144:22]
      InstBoard_1 <= io_WInstNo_1; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_2 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_2) begin // @[RF.scala 144:22]
      InstBoard_2 <= io_WInstNo_2; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_3 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_3) begin // @[RF.scala 144:22]
      InstBoard_3 <= io_WInstNo_3; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_4 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_4) begin // @[RF.scala 144:22]
      InstBoard_4 <= io_WInstNo_4; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_5 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_5) begin // @[RF.scala 144:22]
      InstBoard_5 <= io_WInstNo_5; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_6 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_6) begin // @[RF.scala 144:22]
      InstBoard_6 <= io_WInstNo_6; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_7 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_7) begin // @[RF.scala 144:22]
      InstBoard_7 <= io_WInstNo_7; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_8 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_8) begin // @[RF.scala 144:22]
      InstBoard_8 <= io_WInstNo_8; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_9 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_9) begin // @[RF.scala 144:22]
      InstBoard_9 <= io_WInstNo_9; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_10 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_10) begin // @[RF.scala 144:22]
      InstBoard_10 <= io_WInstNo_10; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_11 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_11) begin // @[RF.scala 144:22]
      InstBoard_11 <= io_WInstNo_11; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_12 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_12) begin // @[RF.scala 144:22]
      InstBoard_12 <= io_WInstNo_12; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_13 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_13) begin // @[RF.scala 144:22]
      InstBoard_13 <= io_WInstNo_13; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_14 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_14) begin // @[RF.scala 144:22]
      InstBoard_14 <= io_WInstNo_14; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_15 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_15) begin // @[RF.scala 144:22]
      InstBoard_15 <= io_WInstNo_15; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_16 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_16) begin // @[RF.scala 144:22]
      InstBoard_16 <= io_WInstNo_16; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_17 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_17) begin // @[RF.scala 144:22]
      InstBoard_17 <= io_WInstNo_17; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_18 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_18) begin // @[RF.scala 144:22]
      InstBoard_18 <= io_WInstNo_18; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_19 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_19) begin // @[RF.scala 144:22]
      InstBoard_19 <= io_WInstNo_19; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_20 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_20) begin // @[RF.scala 144:22]
      InstBoard_20 <= io_WInstNo_20; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_21 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_21) begin // @[RF.scala 144:22]
      InstBoard_21 <= io_WInstNo_21; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_22 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_22) begin // @[RF.scala 144:22]
      InstBoard_22 <= io_WInstNo_22; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_23 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_23) begin // @[RF.scala 144:22]
      InstBoard_23 <= io_WInstNo_23; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_24 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_24) begin // @[RF.scala 144:22]
      InstBoard_24 <= io_WInstNo_24; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_25 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_25) begin // @[RF.scala 144:22]
      InstBoard_25 <= io_WInstNo_25; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_26 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_26) begin // @[RF.scala 144:22]
      InstBoard_26 <= io_WInstNo_26; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_27 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_27) begin // @[RF.scala 144:22]
      InstBoard_27 <= io_WInstNo_27; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_28 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_28) begin // @[RF.scala 144:22]
      InstBoard_28 <= io_WInstNo_28; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_29 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_29) begin // @[RF.scala 144:22]
      InstBoard_29 <= io_WInstNo_29; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_30 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_30) begin // @[RF.scala 144:22]
      InstBoard_30 <= io_WInstNo_30; // @[RF.scala 145:22]
    end
    if (io_flush | reset) begin // @[RF.scala 153:33]
      InstBoard_31 <= 5'h0; // @[RF.scala 139:21]
    end else if (io_Wen_31) begin // @[RF.scala 144:22]
      InstBoard_31 <= io_WInstNo_31; // @[RF.scala 145:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validBoard_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  validBoard_2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  validBoard_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  validBoard_4 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  validBoard_5 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  validBoard_6 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  validBoard_7 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  validBoard_8 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  validBoard_9 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  validBoard_10 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  validBoard_11 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  validBoard_12 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  validBoard_13 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  validBoard_14 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  validBoard_15 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  validBoard_16 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  validBoard_17 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  validBoard_18 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  validBoard_19 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  validBoard_20 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  validBoard_21 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  validBoard_22 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  validBoard_23 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  validBoard_24 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  validBoard_25 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  validBoard_26 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  validBoard_27 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  validBoard_28 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  validBoard_29 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  validBoard_30 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  validBoard_31 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  InstBoard_1 = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  InstBoard_2 = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  InstBoard_3 = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  InstBoard_4 = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  InstBoard_5 = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  InstBoard_6 = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  InstBoard_7 = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  InstBoard_8 = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  InstBoard_9 = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  InstBoard_10 = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  InstBoard_11 = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  InstBoard_12 = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  InstBoard_13 = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  InstBoard_14 = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  InstBoard_15 = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  InstBoard_16 = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  InstBoard_17 = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  InstBoard_18 = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  InstBoard_19 = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  InstBoard_20 = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  InstBoard_21 = _RAND_51[4:0];
  _RAND_52 = {1{`RANDOM}};
  InstBoard_22 = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  InstBoard_23 = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  InstBoard_24 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  InstBoard_25 = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  InstBoard_26 = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  InstBoard_27 = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  InstBoard_28 = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  InstBoard_29 = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  InstBoard_30 = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  InstBoard_31 = _RAND_61[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstQueue(
  input        clock,
  input        reset,
  input  [4:0] io_setnum,
  input  [4:0] io_clearnum,
  output [4:0] io_HeadPtr,
  output [4:0] io_TailPtr,
  output       io_Flag,
  input        io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] HeadPtr; // @[RF.scala 60:24]
  reg [4:0] TailPtr; // @[RF.scala 61:24]
  reg  FlagNow; // @[RF.scala 62:24]
  wire [5:0] _T_2 = io_setnum + HeadPtr; // @[RF.scala 64:29]
  wire [5:0] _T_3 = io_clearnum + TailPtr; // @[RF.scala 65:31]
  wire [5:0] _T_6 = _T_3 - 6'h20; // @[RF.scala 67:29]
  wire [5:0] _GEN_0 = _T_3 >= 6'h20 ? _T_6 : _T_3; // @[RF.scala 66:36 67:15 69:15]
  wire [5:0] _T_361 = _T_2 - 6'h20; // @[RF.scala 83:28]
  wire [5:0] _GEN_97 = _T_2 >= 6'h20 ? _T_361 : _T_2; // @[RF.scala 82:36 83:15 86:15]
  wire [5:0] _GEN_357 = io_flush | reset ? 6'h0 : _GEN_97; // @[RF.scala 109:15 114:33]
  wire [5:0] _GEN_358 = io_flush | reset ? 6'h0 : _GEN_0; // @[RF.scala 110:15 114:33]
  assign io_HeadPtr = HeadPtr; // @[RF.scala 119:13]
  assign io_TailPtr = TailPtr; // @[RF.scala 120:13]
  assign io_Flag = FlagNow; // @[RF.scala 121:13]
  always @(posedge clock) begin
    if (reset) begin // @[RF.scala 60:24]
      HeadPtr <= 5'h0; // @[RF.scala 60:24]
    end else begin
      HeadPtr <= _GEN_357[4:0];
    end
    if (reset) begin // @[RF.scala 61:24]
      TailPtr <= 5'h0; // @[RF.scala 61:24]
    end else begin
      TailPtr <= _GEN_358[4:0];
    end
    if (reset) begin // @[RF.scala 62:24]
      FlagNow <= 1'h0; // @[RF.scala 62:24]
    end else if (io_flush | reset) begin // @[RF.scala 114:33]
      FlagNow <= 1'h0; // @[RF.scala 111:15]
    end else if (_T_2 >= 6'h20) begin // @[RF.scala 82:36]
      FlagNow <= ~FlagNow; // @[RF.scala 84:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  HeadPtr = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  TailPtr = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  FlagNow = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module new_SIMD_ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input  [63:0] io_in_0_bits_cf_runahead_checkpoint_id,
  input  [4:0]  io_in_0_bits_cf_instrType,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [3:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [2:0]  io_in_0_bits_ctrl_funct3,
  input         io_in_0_bits_ctrl_func24,
  input         io_in_0_bits_ctrl_func23,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc3,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input         io_in_0_bits_ctrl_isMou,
  input  [63:0] io_in_0_bits_data_imm,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_cf_instr,
  input  [38:0] io_in_1_bits_cf_pc,
  input  [38:0] io_in_1_bits_cf_pnpc,
  input         io_in_1_bits_cf_exceptionVec_1,
  input         io_in_1_bits_cf_exceptionVec_2,
  input         io_in_1_bits_cf_exceptionVec_12,
  input         io_in_1_bits_cf_intrVec_0,
  input         io_in_1_bits_cf_intrVec_1,
  input         io_in_1_bits_cf_intrVec_2,
  input         io_in_1_bits_cf_intrVec_3,
  input         io_in_1_bits_cf_intrVec_4,
  input         io_in_1_bits_cf_intrVec_5,
  input         io_in_1_bits_cf_intrVec_6,
  input         io_in_1_bits_cf_intrVec_7,
  input         io_in_1_bits_cf_intrVec_8,
  input         io_in_1_bits_cf_intrVec_9,
  input         io_in_1_bits_cf_intrVec_10,
  input         io_in_1_bits_cf_intrVec_11,
  input  [3:0]  io_in_1_bits_cf_brIdx,
  input         io_in_1_bits_cf_crossPageIPFFix,
  input  [63:0] io_in_1_bits_cf_runahead_checkpoint_id,
  input  [4:0]  io_in_1_bits_cf_instrType,
  input         io_in_1_bits_ctrl_src1Type,
  input         io_in_1_bits_ctrl_src2Type,
  input  [3:0]  io_in_1_bits_ctrl_fuType,
  input  [6:0]  io_in_1_bits_ctrl_fuOpType,
  input  [2:0]  io_in_1_bits_ctrl_funct3,
  input         io_in_1_bits_ctrl_func24,
  input         io_in_1_bits_ctrl_func23,
  input  [4:0]  io_in_1_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_1_bits_ctrl_rfSrc2,
  input  [4:0]  io_in_1_bits_ctrl_rfSrc3,
  input         io_in_1_bits_ctrl_rfWen,
  input  [4:0]  io_in_1_bits_ctrl_rfDest,
  input         io_in_1_bits_ctrl_isMou,
  input  [63:0] io_in_1_bits_data_imm,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [63:0] io_out_0_bits_cf_runahead_checkpoint_id,
  output [4:0]  io_out_0_bits_cf_instrType,
  output [3:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [2:0]  io_out_0_bits_ctrl_funct3,
  output        io_out_0_bits_ctrl_func24,
  output        io_out_0_bits_ctrl_func23,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output        io_out_0_bits_ctrl_isBru,
  output        io_out_0_bits_ctrl_isMou,
  output [63:0] io_out_0_bits_data_src1,
  output [63:0] io_out_0_bits_data_src2,
  output [63:0] io_out_0_bits_data_src3,
  output [63:0] io_out_0_bits_data_imm,
  output [4:0]  io_out_0_bits_InstNo,
  output        io_out_0_bits_InstFlag,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [63:0] io_out_1_bits_cf_instr,
  output [38:0] io_out_1_bits_cf_pc,
  output [38:0] io_out_1_bits_cf_pnpc,
  output        io_out_1_bits_cf_exceptionVec_1,
  output        io_out_1_bits_cf_exceptionVec_2,
  output        io_out_1_bits_cf_exceptionVec_12,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  output [3:0]  io_out_1_bits_cf_brIdx,
  output        io_out_1_bits_cf_crossPageIPFFix,
  output [63:0] io_out_1_bits_cf_runahead_checkpoint_id,
  output [4:0]  io_out_1_bits_cf_instrType,
  output [3:0]  io_out_1_bits_ctrl_fuType,
  output [6:0]  io_out_1_bits_ctrl_fuOpType,
  output [2:0]  io_out_1_bits_ctrl_funct3,
  output        io_out_1_bits_ctrl_func24,
  output        io_out_1_bits_ctrl_func23,
  output        io_out_1_bits_ctrl_rfWen,
  output [4:0]  io_out_1_bits_ctrl_rfDest,
  output        io_out_1_bits_ctrl_isBru,
  output        io_out_1_bits_ctrl_isMou,
  output [63:0] io_out_1_bits_data_src1,
  output [63:0] io_out_1_bits_data_src2,
  output [63:0] io_out_1_bits_data_src3,
  output [63:0] io_out_1_bits_data_imm,
  output [4:0]  io_out_1_bits_InstNo,
  output        io_out_1_bits_InstFlag,
  input         io_wb_rfWen_0,
  input         io_wb_rfWen_1,
  input         io_wb_rfWen_2,
  input         io_wb_rfWen_3,
  input         io_wb_rfWen_4,
  input         io_wb_rfWen_5,
  input         io_wb_rfWen_6,
  input         io_wb_rfWen_7,
  input  [4:0]  io_wb_rfDest_0,
  input  [4:0]  io_wb_rfDest_1,
  input  [4:0]  io_wb_rfDest_2,
  input  [4:0]  io_wb_rfDest_3,
  input  [4:0]  io_wb_rfDest_4,
  input  [4:0]  io_wb_rfDest_5,
  input  [4:0]  io_wb_rfDest_6,
  input  [4:0]  io_wb_rfDest_7,
  input  [63:0] io_wb_WriteData_0,
  input  [63:0] io_wb_WriteData_1,
  input  [63:0] io_wb_WriteData_2,
  input  [63:0] io_wb_WriteData_3,
  input  [63:0] io_wb_WriteData_4,
  input  [63:0] io_wb_WriteData_5,
  input  [63:0] io_wb_WriteData_6,
  input  [63:0] io_wb_WriteData_7,
  output [4:0]  io_wb_rfSrc1_0,
  output [4:0]  io_wb_rfSrc1_1,
  output [4:0]  io_wb_rfSrc2_0,
  output [4:0]  io_wb_rfSrc2_1,
  output [4:0]  io_wb_rfSrc3_0,
  output [4:0]  io_wb_rfSrc3_1,
  input  [63:0] io_wb_ReadData1_0,
  input  [63:0] io_wb_ReadData1_1,
  input  [63:0] io_wb_ReadData2_0,
  input  [63:0] io_wb_ReadData2_1,
  input  [63:0] io_wb_ReadData3_0,
  input  [63:0] io_wb_ReadData3_1,
  input  [4:0]  io_wb_InstNo_0,
  input  [4:0]  io_wb_InstNo_1,
  input  [4:0]  io_wb_InstNo_2,
  input  [4:0]  io_wb_InstNo_3,
  input  [4:0]  io_wb_InstNo_4,
  input  [4:0]  io_wb_InstNo_5,
  input  [4:0]  io_wb_InstNo_6,
  input  [4:0]  io_wb_InstNo_7,
  input         io_forward_0_valid,
  input         io_forward_0_wb_rfWen,
  input  [4:0]  io_forward_0_wb_rfDest,
  input  [63:0] io_forward_0_wb_rfData,
  input  [4:0]  io_forward_0_InstNo,
  input         io_forward_1_valid,
  input         io_forward_1_wb_rfWen,
  input  [4:0]  io_forward_1_wb_rfDest,
  input  [63:0] io_forward_1_wb_rfData,
  input  [4:0]  io_forward_1_InstNo,
  input         io_forward_2_valid,
  input         io_forward_2_wb_rfWen,
  input  [4:0]  io_forward_2_wb_rfDest,
  input  [63:0] io_forward_2_wb_rfData,
  input  [4:0]  io_forward_2_InstNo,
  input         io_forward_3_valid,
  input         io_forward_3_wb_rfWen,
  input  [4:0]  io_forward_3_wb_rfDest,
  input  [63:0] io_forward_3_wb_rfData,
  input  [4:0]  io_forward_3_InstNo,
  input         io_forward_4_valid,
  input         io_forward_4_wb_rfWen,
  input  [4:0]  io_forward_4_wb_rfDest,
  input  [63:0] io_forward_4_wb_rfData,
  input  [4:0]  io_forward_4_InstNo,
  input         io_forward_5_valid,
  input         io_forward_5_wb_rfWen,
  input  [4:0]  io_forward_5_wb_rfDest,
  input  [63:0] io_forward_5_wb_rfData,
  input  [4:0]  io_forward_5_InstNo,
  input         io_forward_6_valid,
  input         io_forward_6_wb_rfWen,
  input  [4:0]  io_forward_6_wb_rfDest,
  input  [63:0] io_forward_6_wb_rfData,
  input  [4:0]  io_forward_6_InstNo,
  input         io_forward_7_valid,
  input         io_forward_7_wb_rfWen,
  input  [4:0]  io_forward_7_wb_rfDest,
  input  [63:0] io_forward_7_wb_rfData,
  input  [4:0]  io_forward_7_InstNo,
  input         io_flush,
  input  [4:0]  io_num_enterwbu,
  output [4:0]  io_TailPtr
);
  wire  InstBoard_clock; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_reset; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_1; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_2; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_3; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_4; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_5; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_6; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_7; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_8; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_9; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_10; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_11; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_12; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_13; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_14; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_15; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_16; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_17; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_18; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_19; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_20; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_21; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_22; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_23; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_24; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_25; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_26; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_27; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_28; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_29; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_30; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_Wen_31; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_1; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_2; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_3; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_4; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_5; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_6; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_7; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_8; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_9; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_10; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_11; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_12; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_13; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_14; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_15; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_16; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_17; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_18; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_19; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_20; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_21; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_22; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_23; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_24; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_25; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_26; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_27; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_28; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_29; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_30; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_clear_31; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_1; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_2; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_3; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_4; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_5; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_6; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_7; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_8; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_9; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_10; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_11; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_12; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_13; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_14; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_15; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_16; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_17; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_18; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_19; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_20; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_21; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_22; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_23; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_24; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_25; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_26; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_27; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_28; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_29; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_30; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_WInstNo_31; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_1; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_2; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_3; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_4; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_5; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_6; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_7; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_8; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_9; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_10; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_11; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_12; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_13; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_14; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_15; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_16; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_17; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_18; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_19; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_20; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_21; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_22; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_23; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_24; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_25; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_26; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_27; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_28; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_29; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_30; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_valid_31; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_1; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_2; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_3; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_4; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_5; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_6; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_7; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_8; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_9; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_10; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_11; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_12; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_13; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_14; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_15; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_16; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_17; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_18; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_19; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_20; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_21; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_22; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_23; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_24; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_25; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_26; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_27; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_28; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_29; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_30; // @[SIMD_ISU.scala 163:27]
  wire [4:0] InstBoard_io_RInstNo_31; // @[SIMD_ISU.scala 163:27]
  wire  InstBoard_io_flush; // @[SIMD_ISU.scala 163:27]
  wire  q_clock; // @[SIMD_ISU.scala 164:19]
  wire  q_reset; // @[SIMD_ISU.scala 164:19]
  wire [4:0] q_io_setnum; // @[SIMD_ISU.scala 164:19]
  wire [4:0] q_io_clearnum; // @[SIMD_ISU.scala 164:19]
  wire [4:0] q_io_HeadPtr; // @[SIMD_ISU.scala 164:19]
  wire [4:0] q_io_TailPtr; // @[SIMD_ISU.scala 164:19]
  wire  q_io_Flag; // @[SIMD_ISU.scala 164:19]
  wire  q_io_flush; // @[SIMD_ISU.scala 164:19]
  wire  forwardRfWen_0 = io_forward_0_wb_rfWen & io_forward_0_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_1 = io_forward_1_wb_rfWen & io_forward_1_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_2 = io_forward_2_wb_rfWen & io_forward_2_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_3 = io_forward_3_wb_rfWen & io_forward_3_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_4 = io_forward_4_wb_rfWen & io_forward_4_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_5 = io_forward_5_wb_rfWen & io_forward_5_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_6 = io_forward_6_wb_rfWen & io_forward_6_valid; // @[SIMD_ISU.scala 177:84]
  wire  forwardRfWen_7 = io_forward_7_wb_rfWen & io_forward_7_valid; // @[SIMD_ISU.scala 177:84]
  wire [4:0] _GEN_1 = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_1 : 5'h0; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_2 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_2 : _GEN_1; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_3 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_3 : _GEN_2; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_4 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_4 : _GEN_3; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_5 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_5 : _GEN_4; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_6 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_6 : _GEN_5; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_7 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_7 : _GEN_6; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_8 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_8 : _GEN_7; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_9 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_9 : _GEN_8; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_10 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_10 : _GEN_9; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_11 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_11 : _GEN_10; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_12 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_12 : _GEN_11; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_13 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_13 : _GEN_12; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_14 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_14 : _GEN_13; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_15 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_15 : _GEN_14; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_16 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_16 : _GEN_15; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_17 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_17 : _GEN_16; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_18 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_18 : _GEN_17; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_19 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_19 : _GEN_18; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_20 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_20 : _GEN_19; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_21 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_21 : _GEN_20; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_22 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_22 : _GEN_21; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_23 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_23 : _GEN_22; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_24 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_24 : _GEN_23; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_25 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_25 : _GEN_24; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_26 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_26 : _GEN_25; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_27 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_27 : _GEN_26; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_28 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_28 : _GEN_27; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_29 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_29 : _GEN_28; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_30 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_30 : _GEN_29; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_31 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_31 : _GEN_30; // @[SIMD_ISU.scala 169:{82,82}]
  wire  _T_8 = _GEN_31 == io_forward_0_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_12 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_0_wb_rfDest & forwardRfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_0 = _T_8 & _T_12; // @[SIMD_ISU.scala 178:140]
  wire  _T_14 = _GEN_31 == io_forward_1_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_18 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_1_wb_rfDest & forwardRfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_1 = _T_14 & _T_18; // @[SIMD_ISU.scala 178:140]
  wire  _T_20 = _GEN_31 == io_forward_2_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_24 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_2_wb_rfDest & forwardRfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_2 = _T_20 & _T_24; // @[SIMD_ISU.scala 178:140]
  wire  _T_26 = _GEN_31 == io_forward_3_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_30 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_3_wb_rfDest & forwardRfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_3 = _T_26 & _T_30; // @[SIMD_ISU.scala 178:140]
  wire  _T_32 = _GEN_31 == io_forward_4_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_36 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_4_wb_rfDest & forwardRfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_4 = _T_32 & _T_36; // @[SIMD_ISU.scala 178:140]
  wire  _T_38 = _GEN_31 == io_forward_5_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_42 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_5_wb_rfDest & forwardRfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_5 = _T_38 & _T_42; // @[SIMD_ISU.scala 178:140]
  wire  _T_44 = _GEN_31 == io_forward_6_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_48 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_6_wb_rfDest & forwardRfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_6 = _T_44 & _T_48; // @[SIMD_ISU.scala 178:140]
  wire  _T_50 = _GEN_31 == io_forward_7_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_54 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_7_wb_rfDest & forwardRfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_0_7 = _T_50 & _T_54; // @[SIMD_ISU.scala 178:140]
  wire [4:0] _GEN_33 = 5'h1 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_1 : 5'h0; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_34 = 5'h2 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_2 : _GEN_33; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_35 = 5'h3 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_3 : _GEN_34; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_36 = 5'h4 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_4 : _GEN_35; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_37 = 5'h5 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_5 : _GEN_36; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_38 = 5'h6 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_6 : _GEN_37; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_39 = 5'h7 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_7 : _GEN_38; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_40 = 5'h8 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_8 : _GEN_39; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_41 = 5'h9 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_9 : _GEN_40; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_42 = 5'ha == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_10 : _GEN_41; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_43 = 5'hb == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_11 : _GEN_42; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_44 = 5'hc == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_12 : _GEN_43; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_45 = 5'hd == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_13 : _GEN_44; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_46 = 5'he == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_14 : _GEN_45; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_47 = 5'hf == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_15 : _GEN_46; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_48 = 5'h10 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_16 : _GEN_47; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_49 = 5'h11 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_17 : _GEN_48; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_50 = 5'h12 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_18 : _GEN_49; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_51 = 5'h13 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_19 : _GEN_50; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_52 = 5'h14 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_20 : _GEN_51; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_53 = 5'h15 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_21 : _GEN_52; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_54 = 5'h16 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_22 : _GEN_53; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_55 = 5'h17 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_23 : _GEN_54; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_56 = 5'h18 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_24 : _GEN_55; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_57 = 5'h19 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_25 : _GEN_56; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_58 = 5'h1a == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_26 : _GEN_57; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_59 = 5'h1b == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_27 : _GEN_58; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_60 = 5'h1c == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_28 : _GEN_59; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_61 = 5'h1d == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_29 : _GEN_60; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_62 = 5'h1e == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_30 : _GEN_61; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_63 = 5'h1f == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_RInstNo_31 : _GEN_62; // @[SIMD_ISU.scala 169:{82,82}]
  wire  _T_56 = _GEN_63 == io_forward_0_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_60 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_0_wb_rfDest & forwardRfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_0 = _T_56 & _T_60; // @[SIMD_ISU.scala 178:140]
  wire  _T_62 = _GEN_63 == io_forward_1_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_66 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_1_wb_rfDest & forwardRfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_1 = _T_62 & _T_66; // @[SIMD_ISU.scala 178:140]
  wire  _T_68 = _GEN_63 == io_forward_2_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_72 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_2_wb_rfDest & forwardRfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_2 = _T_68 & _T_72; // @[SIMD_ISU.scala 178:140]
  wire  _T_74 = _GEN_63 == io_forward_3_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_78 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_3_wb_rfDest & forwardRfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_3 = _T_74 & _T_78; // @[SIMD_ISU.scala 178:140]
  wire  _T_80 = _GEN_63 == io_forward_4_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_84 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_4_wb_rfDest & forwardRfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_4 = _T_80 & _T_84; // @[SIMD_ISU.scala 178:140]
  wire  _T_86 = _GEN_63 == io_forward_5_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_90 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_5_wb_rfDest & forwardRfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_5 = _T_86 & _T_90; // @[SIMD_ISU.scala 178:140]
  wire  _T_92 = _GEN_63 == io_forward_6_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_96 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_6_wb_rfDest & forwardRfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_6 = _T_92 & _T_96; // @[SIMD_ISU.scala 178:140]
  wire  _T_98 = _GEN_63 == io_forward_7_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_102 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_forward_7_wb_rfDest & forwardRfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src1DependEX_1_7 = _T_98 & _T_102; // @[SIMD_ISU.scala 178:140]
  wire [4:0] _GEN_65 = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_1 : 5'h0; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_66 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_2 : _GEN_65; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_67 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_3 : _GEN_66; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_68 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_4 : _GEN_67; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_69 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_5 : _GEN_68; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_70 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_6 : _GEN_69; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_71 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_7 : _GEN_70; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_72 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_8 : _GEN_71; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_73 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_9 : _GEN_72; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_74 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_10 : _GEN_73; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_75 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_11 : _GEN_74; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_76 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_12 : _GEN_75; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_77 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_13 : _GEN_76; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_78 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_14 : _GEN_77; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_79 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_15 : _GEN_78; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_80 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_16 : _GEN_79; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_81 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_17 : _GEN_80; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_82 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_18 : _GEN_81; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_83 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_19 : _GEN_82; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_84 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_20 : _GEN_83; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_85 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_21 : _GEN_84; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_86 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_22 : _GEN_85; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_87 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_23 : _GEN_86; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_88 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_24 : _GEN_87; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_89 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_25 : _GEN_88; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_90 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_26 : _GEN_89; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_91 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_27 : _GEN_90; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_92 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_28 : _GEN_91; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_93 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_29 : _GEN_92; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_94 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_30 : _GEN_93; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_95 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_31 : _GEN_94; // @[SIMD_ISU.scala 169:{82,82}]
  wire  _T_104 = _GEN_95 == io_forward_0_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_108 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_0_wb_rfDest & forwardRfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_0 = _T_104 & _T_108; // @[SIMD_ISU.scala 179:140]
  wire  _T_110 = _GEN_95 == io_forward_1_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_114 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_1_wb_rfDest & forwardRfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_1 = _T_110 & _T_114; // @[SIMD_ISU.scala 179:140]
  wire  _T_116 = _GEN_95 == io_forward_2_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_120 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_2_wb_rfDest & forwardRfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_2 = _T_116 & _T_120; // @[SIMD_ISU.scala 179:140]
  wire  _T_122 = _GEN_95 == io_forward_3_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_126 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_3_wb_rfDest & forwardRfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_3 = _T_122 & _T_126; // @[SIMD_ISU.scala 179:140]
  wire  _T_128 = _GEN_95 == io_forward_4_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_132 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_4_wb_rfDest & forwardRfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_4 = _T_128 & _T_132; // @[SIMD_ISU.scala 179:140]
  wire  _T_134 = _GEN_95 == io_forward_5_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_138 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_5_wb_rfDest & forwardRfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_5 = _T_134 & _T_138; // @[SIMD_ISU.scala 179:140]
  wire  _T_140 = _GEN_95 == io_forward_6_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_144 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_6_wb_rfDest & forwardRfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_6 = _T_140 & _T_144; // @[SIMD_ISU.scala 179:140]
  wire  _T_146 = _GEN_95 == io_forward_7_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_150 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_7_wb_rfDest & forwardRfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_0_7 = _T_146 & _T_150; // @[SIMD_ISU.scala 179:140]
  wire [4:0] _GEN_97 = 5'h1 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_1 : 5'h0; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_98 = 5'h2 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_2 : _GEN_97; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_99 = 5'h3 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_3 : _GEN_98; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_100 = 5'h4 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_4 : _GEN_99; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_101 = 5'h5 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_5 : _GEN_100; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_102 = 5'h6 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_6 : _GEN_101; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_103 = 5'h7 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_7 : _GEN_102; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_104 = 5'h8 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_8 : _GEN_103; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_105 = 5'h9 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_9 : _GEN_104; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_106 = 5'ha == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_10 : _GEN_105; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_107 = 5'hb == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_11 : _GEN_106; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_108 = 5'hc == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_12 : _GEN_107; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_109 = 5'hd == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_13 : _GEN_108; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_110 = 5'he == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_14 : _GEN_109; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_111 = 5'hf == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_15 : _GEN_110; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_112 = 5'h10 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_16 : _GEN_111; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_113 = 5'h11 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_17 : _GEN_112; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_114 = 5'h12 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_18 : _GEN_113; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_115 = 5'h13 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_19 : _GEN_114; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_116 = 5'h14 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_20 : _GEN_115; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_117 = 5'h15 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_21 : _GEN_116; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_118 = 5'h16 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_22 : _GEN_117; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_119 = 5'h17 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_23 : _GEN_118; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_120 = 5'h18 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_24 : _GEN_119; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_121 = 5'h19 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_25 : _GEN_120; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_122 = 5'h1a == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_26 : _GEN_121; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_123 = 5'h1b == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_27 : _GEN_122; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_124 = 5'h1c == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_28 : _GEN_123; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_125 = 5'h1d == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_29 : _GEN_124; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_126 = 5'h1e == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_30 : _GEN_125; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_127 = 5'h1f == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_RInstNo_31 : _GEN_126; // @[SIMD_ISU.scala 169:{82,82}]
  wire  _T_152 = _GEN_127 == io_forward_0_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_156 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_0_wb_rfDest & forwardRfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_0 = _T_152 & _T_156; // @[SIMD_ISU.scala 179:140]
  wire  _T_158 = _GEN_127 == io_forward_1_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_162 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_1_wb_rfDest & forwardRfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_1 = _T_158 & _T_162; // @[SIMD_ISU.scala 179:140]
  wire  _T_164 = _GEN_127 == io_forward_2_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_168 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_2_wb_rfDest & forwardRfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_2 = _T_164 & _T_168; // @[SIMD_ISU.scala 179:140]
  wire  _T_170 = _GEN_127 == io_forward_3_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_174 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_3_wb_rfDest & forwardRfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_3 = _T_170 & _T_174; // @[SIMD_ISU.scala 179:140]
  wire  _T_176 = _GEN_127 == io_forward_4_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_180 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_4_wb_rfDest & forwardRfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_4 = _T_176 & _T_180; // @[SIMD_ISU.scala 179:140]
  wire  _T_182 = _GEN_127 == io_forward_5_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_186 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_5_wb_rfDest & forwardRfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_5 = _T_182 & _T_186; // @[SIMD_ISU.scala 179:140]
  wire  _T_188 = _GEN_127 == io_forward_6_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_192 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_6_wb_rfDest & forwardRfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_6 = _T_188 & _T_192; // @[SIMD_ISU.scala 179:140]
  wire  _T_194 = _GEN_127 == io_forward_7_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_198 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_forward_7_wb_rfDest & forwardRfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src2DependEX_1_7 = _T_194 & _T_198; // @[SIMD_ISU.scala 179:140]
  wire  _T_200 = _GEN_31 == io_wb_InstNo_0; // @[SIMD_ISU.scala 169:82]
  wire  _T_204 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_0 & io_wb_rfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_0 = _T_200 & _T_204; // @[SIMD_ISU.scala 180:135]
  wire  _T_206 = _GEN_31 == io_wb_InstNo_1; // @[SIMD_ISU.scala 169:82]
  wire  _T_210 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_1 & io_wb_rfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_1 = _T_206 & _T_210; // @[SIMD_ISU.scala 180:135]
  wire  _T_212 = _GEN_31 == io_wb_InstNo_2; // @[SIMD_ISU.scala 169:82]
  wire  _T_216 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_2 & io_wb_rfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_2 = _T_212 & _T_216; // @[SIMD_ISU.scala 180:135]
  wire  _T_218 = _GEN_31 == io_wb_InstNo_3; // @[SIMD_ISU.scala 169:82]
  wire  _T_222 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_3 & io_wb_rfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_3 = _T_218 & _T_222; // @[SIMD_ISU.scala 180:135]
  wire  _T_224 = _GEN_31 == io_wb_InstNo_4; // @[SIMD_ISU.scala 169:82]
  wire  _T_228 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_4 & io_wb_rfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_4 = _T_224 & _T_228; // @[SIMD_ISU.scala 180:135]
  wire  _T_230 = _GEN_31 == io_wb_InstNo_5; // @[SIMD_ISU.scala 169:82]
  wire  _T_234 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_5 & io_wb_rfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_5 = _T_230 & _T_234; // @[SIMD_ISU.scala 180:135]
  wire  _T_236 = _GEN_31 == io_wb_InstNo_6; // @[SIMD_ISU.scala 169:82]
  wire  _T_240 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_6 & io_wb_rfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_6 = _T_236 & _T_240; // @[SIMD_ISU.scala 180:135]
  wire  _T_242 = _GEN_31 == io_wb_InstNo_7; // @[SIMD_ISU.scala 169:82]
  wire  _T_246 = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest_7 & io_wb_rfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_0_7 = _T_242 & _T_246; // @[SIMD_ISU.scala 180:135]
  wire  _T_248 = _GEN_63 == io_wb_InstNo_0; // @[SIMD_ISU.scala 169:82]
  wire  _T_252 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_0 & io_wb_rfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_0 = _T_248 & _T_252; // @[SIMD_ISU.scala 180:135]
  wire  _T_254 = _GEN_63 == io_wb_InstNo_1; // @[SIMD_ISU.scala 169:82]
  wire  _T_258 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_1 & io_wb_rfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_1 = _T_254 & _T_258; // @[SIMD_ISU.scala 180:135]
  wire  _T_260 = _GEN_63 == io_wb_InstNo_2; // @[SIMD_ISU.scala 169:82]
  wire  _T_264 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_2 & io_wb_rfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_2 = _T_260 & _T_264; // @[SIMD_ISU.scala 180:135]
  wire  _T_266 = _GEN_63 == io_wb_InstNo_3; // @[SIMD_ISU.scala 169:82]
  wire  _T_270 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_3 & io_wb_rfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_3 = _T_266 & _T_270; // @[SIMD_ISU.scala 180:135]
  wire  _T_272 = _GEN_63 == io_wb_InstNo_4; // @[SIMD_ISU.scala 169:82]
  wire  _T_276 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_4 & io_wb_rfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_4 = _T_272 & _T_276; // @[SIMD_ISU.scala 180:135]
  wire  _T_278 = _GEN_63 == io_wb_InstNo_5; // @[SIMD_ISU.scala 169:82]
  wire  _T_282 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_5 & io_wb_rfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_5 = _T_278 & _T_282; // @[SIMD_ISU.scala 180:135]
  wire  _T_284 = _GEN_63 == io_wb_InstNo_6; // @[SIMD_ISU.scala 169:82]
  wire  _T_288 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_6 & io_wb_rfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_6 = _T_284 & _T_288; // @[SIMD_ISU.scala 180:135]
  wire  _T_290 = _GEN_63 == io_wb_InstNo_7; // @[SIMD_ISU.scala 169:82]
  wire  _T_294 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_wb_rfDest_7 & io_wb_rfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src1DependWB_1_7 = _T_290 & _T_294; // @[SIMD_ISU.scala 180:135]
  wire  _T_296 = _GEN_95 == io_wb_InstNo_0; // @[SIMD_ISU.scala 169:82]
  wire  _T_300 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_0 & io_wb_rfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_0 = _T_296 & _T_300; // @[SIMD_ISU.scala 181:135]
  wire  _T_302 = _GEN_95 == io_wb_InstNo_1; // @[SIMD_ISU.scala 169:82]
  wire  _T_306 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_1 & io_wb_rfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_1 = _T_302 & _T_306; // @[SIMD_ISU.scala 181:135]
  wire  _T_308 = _GEN_95 == io_wb_InstNo_2; // @[SIMD_ISU.scala 169:82]
  wire  _T_312 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_2 & io_wb_rfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_2 = _T_308 & _T_312; // @[SIMD_ISU.scala 181:135]
  wire  _T_314 = _GEN_95 == io_wb_InstNo_3; // @[SIMD_ISU.scala 169:82]
  wire  _T_318 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_3 & io_wb_rfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_3 = _T_314 & _T_318; // @[SIMD_ISU.scala 181:135]
  wire  _T_320 = _GEN_95 == io_wb_InstNo_4; // @[SIMD_ISU.scala 169:82]
  wire  _T_324 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_4 & io_wb_rfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_4 = _T_320 & _T_324; // @[SIMD_ISU.scala 181:135]
  wire  _T_326 = _GEN_95 == io_wb_InstNo_5; // @[SIMD_ISU.scala 169:82]
  wire  _T_330 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_5 & io_wb_rfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_5 = _T_326 & _T_330; // @[SIMD_ISU.scala 181:135]
  wire  _T_332 = _GEN_95 == io_wb_InstNo_6; // @[SIMD_ISU.scala 169:82]
  wire  _T_336 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_6 & io_wb_rfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_6 = _T_332 & _T_336; // @[SIMD_ISU.scala 181:135]
  wire  _T_338 = _GEN_95 == io_wb_InstNo_7; // @[SIMD_ISU.scala 169:82]
  wire  _T_342 = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest_7 & io_wb_rfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_0_7 = _T_338 & _T_342; // @[SIMD_ISU.scala 181:135]
  wire  _T_344 = _GEN_127 == io_wb_InstNo_0; // @[SIMD_ISU.scala 169:82]
  wire  _T_348 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_0 & io_wb_rfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_0 = _T_344 & _T_348; // @[SIMD_ISU.scala 181:135]
  wire  _T_350 = _GEN_127 == io_wb_InstNo_1; // @[SIMD_ISU.scala 169:82]
  wire  _T_354 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_1 & io_wb_rfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_1 = _T_350 & _T_354; // @[SIMD_ISU.scala 181:135]
  wire  _T_356 = _GEN_127 == io_wb_InstNo_2; // @[SIMD_ISU.scala 169:82]
  wire  _T_360 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_2 & io_wb_rfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_2 = _T_356 & _T_360; // @[SIMD_ISU.scala 181:135]
  wire  _T_362 = _GEN_127 == io_wb_InstNo_3; // @[SIMD_ISU.scala 169:82]
  wire  _T_366 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_3 & io_wb_rfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_3 = _T_362 & _T_366; // @[SIMD_ISU.scala 181:135]
  wire  _T_368 = _GEN_127 == io_wb_InstNo_4; // @[SIMD_ISU.scala 169:82]
  wire  _T_372 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_4 & io_wb_rfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_4 = _T_368 & _T_372; // @[SIMD_ISU.scala 181:135]
  wire  _T_374 = _GEN_127 == io_wb_InstNo_5; // @[SIMD_ISU.scala 169:82]
  wire  _T_378 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_5 & io_wb_rfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_5 = _T_374 & _T_378; // @[SIMD_ISU.scala 181:135]
  wire  _T_380 = _GEN_127 == io_wb_InstNo_6; // @[SIMD_ISU.scala 169:82]
  wire  _T_384 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_6 & io_wb_rfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_6 = _T_380 & _T_384; // @[SIMD_ISU.scala 181:135]
  wire  _T_386 = _GEN_127 == io_wb_InstNo_7; // @[SIMD_ISU.scala 169:82]
  wire  _T_390 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_wb_rfDest_7 & io_wb_rfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  src2DependWB_1_7 = _T_386 & _T_390; // @[SIMD_ISU.scala 181:135]
  wire  _GEN_130 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_2 : 5'h1 == io_in_0_bits_ctrl_rfSrc1 &
    InstBoard_io_valid_1; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_131 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_3 : _GEN_130; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_132 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_4 : _GEN_131; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_133 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_5 : _GEN_132; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_134 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_6 : _GEN_133; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_135 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_7 : _GEN_134; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_136 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_8 : _GEN_135; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_137 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_9 : _GEN_136; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_138 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_10 : _GEN_137; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_139 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_11 : _GEN_138; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_140 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_12 : _GEN_139; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_141 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_13 : _GEN_140; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_142 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_14 : _GEN_141; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_143 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_15 : _GEN_142; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_144 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_16 : _GEN_143; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_145 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_17 : _GEN_144; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_146 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_18 : _GEN_145; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_147 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_19 : _GEN_146; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_148 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_20 : _GEN_147; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_149 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_21 : _GEN_148; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_150 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_22 : _GEN_149; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_151 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_23 : _GEN_150; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_152 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_24 : _GEN_151; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_153 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_25 : _GEN_152; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_154 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_26 : _GEN_153; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_155 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_27 : _GEN_154; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_156 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_28 : _GEN_155; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_157 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_29 : _GEN_156; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_158 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_30 : _GEN_157; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_159 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? InstBoard_io_valid_31 : _GEN_158; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _T_399 = src1DependEX_0_0 | src1DependEX_0_1 | src1DependEX_0_2 | src1DependEX_0_3 | src1DependEX_0_4 |
    src1DependEX_0_5 | src1DependEX_0_6 | src1DependEX_0_7; // @[SIMD_ISU.scala 183:113]
  wire  _T_407 = src1DependWB_0_0 | src1DependWB_0_1 | src1DependWB_0_2 | src1DependWB_0_3 | src1DependWB_0_4 |
    src1DependWB_0_5 | src1DependWB_0_6 | src1DependWB_0_7; // @[SIMD_ISU.scala 183:143]
  wire  src1Ready_0 = ~_GEN_159 | (src1DependEX_0_0 | src1DependEX_0_1 | src1DependEX_0_2 | src1DependEX_0_3 |
    src1DependEX_0_4 | src1DependEX_0_5 | src1DependEX_0_6 | src1DependEX_0_7) | (src1DependWB_0_0 | src1DependWB_0_1 |
    src1DependWB_0_2 | src1DependWB_0_3 | src1DependWB_0_4 | src1DependWB_0_5 | src1DependWB_0_6 | src1DependWB_0_7); // @[SIMD_ISU.scala 183:117]
  wire  _GEN_162 = 5'h2 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_2 : 5'h1 == io_in_1_bits_ctrl_rfSrc1 &
    InstBoard_io_valid_1; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_163 = 5'h3 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_3 : _GEN_162; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_164 = 5'h4 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_4 : _GEN_163; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_165 = 5'h5 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_5 : _GEN_164; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_166 = 5'h6 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_6 : _GEN_165; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_167 = 5'h7 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_7 : _GEN_166; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_168 = 5'h8 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_8 : _GEN_167; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_169 = 5'h9 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_9 : _GEN_168; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_170 = 5'ha == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_10 : _GEN_169; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_171 = 5'hb == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_11 : _GEN_170; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_172 = 5'hc == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_12 : _GEN_171; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_173 = 5'hd == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_13 : _GEN_172; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_174 = 5'he == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_14 : _GEN_173; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_175 = 5'hf == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_15 : _GEN_174; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_176 = 5'h10 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_16 : _GEN_175; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_177 = 5'h11 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_17 : _GEN_176; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_178 = 5'h12 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_18 : _GEN_177; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_179 = 5'h13 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_19 : _GEN_178; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_180 = 5'h14 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_20 : _GEN_179; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_181 = 5'h15 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_21 : _GEN_180; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_182 = 5'h16 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_22 : _GEN_181; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_183 = 5'h17 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_23 : _GEN_182; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_184 = 5'h18 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_24 : _GEN_183; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_185 = 5'h19 == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_25 : _GEN_184; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_186 = 5'h1a == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_26 : _GEN_185; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_187 = 5'h1b == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_27 : _GEN_186; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_188 = 5'h1c == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_28 : _GEN_187; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_189 = 5'h1d == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_29 : _GEN_188; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_190 = 5'h1e == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_30 : _GEN_189; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _GEN_191 = 5'h1f == io_in_1_bits_ctrl_rfSrc1 ? InstBoard_io_valid_31 : _GEN_190; // @[SIMD_ISU.scala 183:{57,57}]
  wire  _T_416 = src1DependEX_1_0 | src1DependEX_1_1 | src1DependEX_1_2 | src1DependEX_1_3 | src1DependEX_1_4 |
    src1DependEX_1_5 | src1DependEX_1_6 | src1DependEX_1_7; // @[SIMD_ISU.scala 183:113]
  wire  _T_424 = src1DependWB_1_0 | src1DependWB_1_1 | src1DependWB_1_2 | src1DependWB_1_3 | src1DependWB_1_4 |
    src1DependWB_1_5 | src1DependWB_1_6 | src1DependWB_1_7; // @[SIMD_ISU.scala 183:143]
  wire  src1Ready_1 = ~_GEN_191 | (src1DependEX_1_0 | src1DependEX_1_1 | src1DependEX_1_2 | src1DependEX_1_3 |
    src1DependEX_1_4 | src1DependEX_1_5 | src1DependEX_1_6 | src1DependEX_1_7) | (src1DependWB_1_0 | src1DependWB_1_1 |
    src1DependWB_1_2 | src1DependWB_1_3 | src1DependWB_1_4 | src1DependWB_1_5 | src1DependWB_1_6 | src1DependWB_1_7); // @[SIMD_ISU.scala 183:117]
  wire  _GEN_194 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_2 : 5'h1 == io_in_0_bits_ctrl_rfSrc2 &
    InstBoard_io_valid_1; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_195 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_3 : _GEN_194; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_196 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_4 : _GEN_195; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_197 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_5 : _GEN_196; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_198 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_6 : _GEN_197; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_199 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_7 : _GEN_198; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_200 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_8 : _GEN_199; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_201 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_9 : _GEN_200; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_202 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_10 : _GEN_201; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_203 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_11 : _GEN_202; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_204 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_12 : _GEN_203; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_205 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_13 : _GEN_204; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_206 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_14 : _GEN_205; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_207 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_15 : _GEN_206; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_208 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_16 : _GEN_207; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_209 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_17 : _GEN_208; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_210 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_18 : _GEN_209; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_211 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_19 : _GEN_210; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_212 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_20 : _GEN_211; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_213 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_21 : _GEN_212; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_214 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_22 : _GEN_213; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_215 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_23 : _GEN_214; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_216 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_24 : _GEN_215; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_217 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_25 : _GEN_216; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_218 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_26 : _GEN_217; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_219 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_27 : _GEN_218; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_220 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_28 : _GEN_219; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_221 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_29 : _GEN_220; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_222 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_30 : _GEN_221; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_223 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? InstBoard_io_valid_31 : _GEN_222; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _T_433 = src2DependEX_0_0 | src2DependEX_0_1 | src2DependEX_0_2 | src2DependEX_0_3 | src2DependEX_0_4 |
    src2DependEX_0_5 | src2DependEX_0_6 | src2DependEX_0_7; // @[SIMD_ISU.scala 184:113]
  wire  _T_441 = src2DependWB_0_0 | src2DependWB_0_1 | src2DependWB_0_2 | src2DependWB_0_3 | src2DependWB_0_4 |
    src2DependWB_0_5 | src2DependWB_0_6 | src2DependWB_0_7; // @[SIMD_ISU.scala 184:143]
  wire  src2Ready_0 = ~_GEN_223 | (src2DependEX_0_0 | src2DependEX_0_1 | src2DependEX_0_2 | src2DependEX_0_3 |
    src2DependEX_0_4 | src2DependEX_0_5 | src2DependEX_0_6 | src2DependEX_0_7) | (src2DependWB_0_0 | src2DependWB_0_1 |
    src2DependWB_0_2 | src2DependWB_0_3 | src2DependWB_0_4 | src2DependWB_0_5 | src2DependWB_0_6 | src2DependWB_0_7); // @[SIMD_ISU.scala 184:117]
  wire  _GEN_226 = 5'h2 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_2 : 5'h1 == io_in_1_bits_ctrl_rfSrc2 &
    InstBoard_io_valid_1; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_227 = 5'h3 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_3 : _GEN_226; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_228 = 5'h4 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_4 : _GEN_227; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_229 = 5'h5 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_5 : _GEN_228; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_230 = 5'h6 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_6 : _GEN_229; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_231 = 5'h7 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_7 : _GEN_230; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_232 = 5'h8 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_8 : _GEN_231; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_233 = 5'h9 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_9 : _GEN_232; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_234 = 5'ha == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_10 : _GEN_233; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_235 = 5'hb == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_11 : _GEN_234; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_236 = 5'hc == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_12 : _GEN_235; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_237 = 5'hd == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_13 : _GEN_236; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_238 = 5'he == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_14 : _GEN_237; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_239 = 5'hf == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_15 : _GEN_238; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_240 = 5'h10 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_16 : _GEN_239; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_241 = 5'h11 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_17 : _GEN_240; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_242 = 5'h12 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_18 : _GEN_241; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_243 = 5'h13 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_19 : _GEN_242; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_244 = 5'h14 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_20 : _GEN_243; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_245 = 5'h15 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_21 : _GEN_244; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_246 = 5'h16 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_22 : _GEN_245; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_247 = 5'h17 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_23 : _GEN_246; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_248 = 5'h18 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_24 : _GEN_247; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_249 = 5'h19 == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_25 : _GEN_248; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_250 = 5'h1a == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_26 : _GEN_249; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_251 = 5'h1b == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_27 : _GEN_250; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_252 = 5'h1c == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_28 : _GEN_251; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_253 = 5'h1d == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_29 : _GEN_252; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_254 = 5'h1e == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_30 : _GEN_253; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _GEN_255 = 5'h1f == io_in_1_bits_ctrl_rfSrc2 ? InstBoard_io_valid_31 : _GEN_254; // @[SIMD_ISU.scala 184:{57,57}]
  wire  _T_450 = src2DependEX_1_0 | src2DependEX_1_1 | src2DependEX_1_2 | src2DependEX_1_3 | src2DependEX_1_4 |
    src2DependEX_1_5 | src2DependEX_1_6 | src2DependEX_1_7; // @[SIMD_ISU.scala 184:113]
  wire  _T_458 = src2DependWB_1_0 | src2DependWB_1_1 | src2DependWB_1_2 | src2DependWB_1_3 | src2DependWB_1_4 |
    src2DependWB_1_5 | src2DependWB_1_6 | src2DependWB_1_7; // @[SIMD_ISU.scala 184:143]
  wire  src2Ready_1 = ~_GEN_255 | (src2DependEX_1_0 | src2DependEX_1_1 | src2DependEX_1_2 | src2DependEX_1_3 |
    src2DependEX_1_4 | src2DependEX_1_5 | src2DependEX_1_6 | src2DependEX_1_7) | (src2DependWB_1_0 | src2DependWB_1_1 |
    src2DependWB_1_2 | src2DependWB_1_3 | src2DependWB_1_4 | src2DependWB_1_5 | src2DependWB_1_6 | src2DependWB_1_7); // @[SIMD_ISU.scala 184:117]
  wire  _T_464 = io_in_1_bits_ctrl_rfSrc1 != 5'h0 & io_in_1_bits_ctrl_rfSrc1 == io_in_0_bits_ctrl_rfDest &
    io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 166:102]
  wire  _T_468 = io_in_1_bits_ctrl_rfSrc2 != 5'h0 & io_in_1_bits_ctrl_rfSrc2 == io_in_0_bits_ctrl_rfDest &
    io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 166:102]
  wire  _T_473 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_in_0_bits_ctrl_rfDest &
    io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 166:102]
  wire  RAWinIssue_1 = io_in_0_valid & (_T_464 | _T_468 | _T_473); // @[SIMD_ISU.scala 189:90]
  wire  _T_480 = io_in_0_bits_ctrl_fuType == 4'h1 | io_in_0_bits_ctrl_fuType == 4'h8; // @[SIMD_ISU.scala 198:135]
  wire  FrontHasCsrMouOp_1 = io_in_0_valid & (io_in_0_bits_ctrl_fuType == 4'h1 | io_in_0_bits_ctrl_fuType == 4'h8); // @[SIMD_ISU.scala 198:90]
  wire  FrontisClear_1 = ~io_in_0_valid; // @[SIMD_ISU.scala 206:75]
  wire  _GEN_386 = 5'h2 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_2 : 5'h1 == io_in_0_bits_ctrl_rfSrc3 &
    InstBoard_io_valid_1; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_387 = 5'h3 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_3 : _GEN_386; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_388 = 5'h4 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_4 : _GEN_387; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_389 = 5'h5 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_5 : _GEN_388; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_390 = 5'h6 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_6 : _GEN_389; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_391 = 5'h7 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_7 : _GEN_390; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_392 = 5'h8 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_8 : _GEN_391; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_393 = 5'h9 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_9 : _GEN_392; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_394 = 5'ha == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_10 : _GEN_393; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_395 = 5'hb == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_11 : _GEN_394; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_396 = 5'hc == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_12 : _GEN_395; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_397 = 5'hd == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_13 : _GEN_396; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_398 = 5'he == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_14 : _GEN_397; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_399 = 5'hf == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_15 : _GEN_398; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_400 = 5'h10 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_16 : _GEN_399; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_401 = 5'h11 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_17 : _GEN_400; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_402 = 5'h12 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_18 : _GEN_401; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_403 = 5'h13 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_19 : _GEN_402; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_404 = 5'h14 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_20 : _GEN_403; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_405 = 5'h15 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_21 : _GEN_404; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_406 = 5'h16 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_22 : _GEN_405; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_407 = 5'h17 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_23 : _GEN_406; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_408 = 5'h18 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_24 : _GEN_407; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_409 = 5'h19 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_25 : _GEN_408; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_410 = 5'h1a == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_26 : _GEN_409; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_411 = 5'h1b == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_27 : _GEN_410; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_412 = 5'h1c == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_28 : _GEN_411; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_413 = 5'h1d == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_29 : _GEN_412; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_414 = 5'h1e == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_30 : _GEN_413; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_415 = 5'h1f == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_valid_31 : _GEN_414; // @[SIMD_ISU.scala 261:{49,49}]
  wire [4:0] _GEN_321 = 5'h1 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_1 : 5'h0; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_322 = 5'h2 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_2 : _GEN_321; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_323 = 5'h3 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_3 : _GEN_322; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_324 = 5'h4 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_4 : _GEN_323; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_325 = 5'h5 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_5 : _GEN_324; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_326 = 5'h6 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_6 : _GEN_325; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_327 = 5'h7 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_7 : _GEN_326; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_328 = 5'h8 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_8 : _GEN_327; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_329 = 5'h9 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_9 : _GEN_328; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_330 = 5'ha == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_10 : _GEN_329; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_331 = 5'hb == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_11 : _GEN_330; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_332 = 5'hc == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_12 : _GEN_331; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_333 = 5'hd == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_13 : _GEN_332; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_334 = 5'he == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_14 : _GEN_333; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_335 = 5'hf == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_15 : _GEN_334; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_336 = 5'h10 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_16 : _GEN_335; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_337 = 5'h11 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_17 : _GEN_336; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_338 = 5'h12 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_18 : _GEN_337; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_339 = 5'h13 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_19 : _GEN_338; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_340 = 5'h14 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_20 : _GEN_339; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_341 = 5'h15 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_21 : _GEN_340; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_342 = 5'h16 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_22 : _GEN_341; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_343 = 5'h17 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_23 : _GEN_342; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_344 = 5'h18 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_24 : _GEN_343; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_345 = 5'h19 == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_25 : _GEN_344; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_346 = 5'h1a == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_26 : _GEN_345; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_347 = 5'h1b == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_27 : _GEN_346; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_348 = 5'h1c == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_28 : _GEN_347; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_349 = 5'h1d == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_29 : _GEN_348; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_350 = 5'h1e == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_30 : _GEN_349; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_351 = 5'h1f == io_in_0_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_31 : _GEN_350; // @[SIMD_ISU.scala 169:{82,82}]
  wire  _T_820 = _GEN_351 == io_forward_0_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_824 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_0_wb_rfDest & forwardRfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  _T_825 = _T_820 & _T_824; // @[SIMD_ISU.scala 259:140]
  wire  _T_826 = _GEN_351 == io_forward_1_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_830 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_1_wb_rfDest & forwardRfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  _T_831 = _T_826 & _T_830; // @[SIMD_ISU.scala 259:140]
  wire  _T_832 = _GEN_351 == io_forward_2_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_836 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_2_wb_rfDest & forwardRfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  _T_837 = _T_832 & _T_836; // @[SIMD_ISU.scala 259:140]
  wire  _T_838 = _GEN_351 == io_forward_3_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_842 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_3_wb_rfDest & forwardRfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  _T_843 = _T_838 & _T_842; // @[SIMD_ISU.scala 259:140]
  wire  _T_844 = _GEN_351 == io_forward_4_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_848 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_4_wb_rfDest & forwardRfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  _T_849 = _T_844 & _T_848; // @[SIMD_ISU.scala 259:140]
  wire  _T_850 = _GEN_351 == io_forward_5_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_854 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_5_wb_rfDest & forwardRfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  _T_855 = _T_850 & _T_854; // @[SIMD_ISU.scala 259:140]
  wire  _T_856 = _GEN_351 == io_forward_6_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_860 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_6_wb_rfDest & forwardRfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  _T_861 = _T_856 & _T_860; // @[SIMD_ISU.scala 259:140]
  wire  _T_862 = _GEN_351 == io_forward_7_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_866 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_forward_7_wb_rfDest & forwardRfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  _T_867 = _T_862 & _T_866; // @[SIMD_ISU.scala 259:140]
  wire  _T_1019 = _T_825 | _T_831 | _T_837 | _T_843 | _T_849 | _T_855 | _T_861 | _T_867; // @[SIMD_ISU.scala 261:105]
  wire  _T_916 = _GEN_351 == io_wb_InstNo_0; // @[SIMD_ISU.scala 169:82]
  wire  _T_920 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_0 & io_wb_rfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  _T_921 = _T_916 & _T_920; // @[SIMD_ISU.scala 260:135]
  wire  _T_922 = _GEN_351 == io_wb_InstNo_1; // @[SIMD_ISU.scala 169:82]
  wire  _T_926 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_1 & io_wb_rfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  _T_927 = _T_922 & _T_926; // @[SIMD_ISU.scala 260:135]
  wire  _T_928 = _GEN_351 == io_wb_InstNo_2; // @[SIMD_ISU.scala 169:82]
  wire  _T_932 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_2 & io_wb_rfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  _T_933 = _T_928 & _T_932; // @[SIMD_ISU.scala 260:135]
  wire  _T_934 = _GEN_351 == io_wb_InstNo_3; // @[SIMD_ISU.scala 169:82]
  wire  _T_938 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_3 & io_wb_rfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  _T_939 = _T_934 & _T_938; // @[SIMD_ISU.scala 260:135]
  wire  _T_940 = _GEN_351 == io_wb_InstNo_4; // @[SIMD_ISU.scala 169:82]
  wire  _T_944 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_4 & io_wb_rfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  _T_945 = _T_940 & _T_944; // @[SIMD_ISU.scala 260:135]
  wire  _T_946 = _GEN_351 == io_wb_InstNo_5; // @[SIMD_ISU.scala 169:82]
  wire  _T_950 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_5 & io_wb_rfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  _T_951 = _T_946 & _T_950; // @[SIMD_ISU.scala 260:135]
  wire  _T_952 = _GEN_351 == io_wb_InstNo_6; // @[SIMD_ISU.scala 169:82]
  wire  _T_956 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_6 & io_wb_rfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  _T_957 = _T_952 & _T_956; // @[SIMD_ISU.scala 260:135]
  wire  _T_958 = _GEN_351 == io_wb_InstNo_7; // @[SIMD_ISU.scala 169:82]
  wire  _T_962 = io_in_0_bits_ctrl_rfSrc3 != 5'h0 & io_in_0_bits_ctrl_rfSrc3 == io_wb_rfDest_7 & io_wb_rfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  _T_963 = _T_958 & _T_962; // @[SIMD_ISU.scala 260:135]
  wire  _T_1027 = _T_921 | _T_927 | _T_933 | _T_939 | _T_945 | _T_951 | _T_957 | _T_963; // @[SIMD_ISU.scala 261:135]
  wire  src3Ready_0 = ~_GEN_415 | (_T_825 | _T_831 | _T_837 | _T_843 | _T_849 | _T_855 | _T_861 | _T_867) | (_T_921 |
    _T_927 | _T_933 | _T_939 | _T_945 | _T_951 | _T_957 | _T_963); // @[SIMD_ISU.scala 261:109]
  wire  _GEN_418 = 5'h2 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_2 : 5'h1 == io_in_1_bits_ctrl_rfSrc3 &
    InstBoard_io_valid_1; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_419 = 5'h3 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_3 : _GEN_418; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_420 = 5'h4 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_4 : _GEN_419; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_421 = 5'h5 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_5 : _GEN_420; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_422 = 5'h6 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_6 : _GEN_421; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_423 = 5'h7 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_7 : _GEN_422; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_424 = 5'h8 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_8 : _GEN_423; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_425 = 5'h9 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_9 : _GEN_424; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_426 = 5'ha == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_10 : _GEN_425; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_427 = 5'hb == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_11 : _GEN_426; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_428 = 5'hc == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_12 : _GEN_427; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_429 = 5'hd == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_13 : _GEN_428; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_430 = 5'he == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_14 : _GEN_429; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_431 = 5'hf == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_15 : _GEN_430; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_432 = 5'h10 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_16 : _GEN_431; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_433 = 5'h11 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_17 : _GEN_432; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_434 = 5'h12 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_18 : _GEN_433; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_435 = 5'h13 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_19 : _GEN_434; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_436 = 5'h14 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_20 : _GEN_435; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_437 = 5'h15 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_21 : _GEN_436; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_438 = 5'h16 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_22 : _GEN_437; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_439 = 5'h17 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_23 : _GEN_438; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_440 = 5'h18 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_24 : _GEN_439; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_441 = 5'h19 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_25 : _GEN_440; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_442 = 5'h1a == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_26 : _GEN_441; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_443 = 5'h1b == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_27 : _GEN_442; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_444 = 5'h1c == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_28 : _GEN_443; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_445 = 5'h1d == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_29 : _GEN_444; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_446 = 5'h1e == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_30 : _GEN_445; // @[SIMD_ISU.scala 261:{49,49}]
  wire  _GEN_447 = 5'h1f == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_valid_31 : _GEN_446; // @[SIMD_ISU.scala 261:{49,49}]
  wire [4:0] _GEN_353 = 5'h1 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_1 : 5'h0; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_354 = 5'h2 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_2 : _GEN_353; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_355 = 5'h3 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_3 : _GEN_354; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_356 = 5'h4 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_4 : _GEN_355; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_357 = 5'h5 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_5 : _GEN_356; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_358 = 5'h6 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_6 : _GEN_357; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_359 = 5'h7 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_7 : _GEN_358; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_360 = 5'h8 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_8 : _GEN_359; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_361 = 5'h9 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_9 : _GEN_360; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_362 = 5'ha == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_10 : _GEN_361; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_363 = 5'hb == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_11 : _GEN_362; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_364 = 5'hc == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_12 : _GEN_363; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_365 = 5'hd == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_13 : _GEN_364; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_366 = 5'he == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_14 : _GEN_365; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_367 = 5'hf == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_15 : _GEN_366; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_368 = 5'h10 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_16 : _GEN_367; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_369 = 5'h11 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_17 : _GEN_368; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_370 = 5'h12 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_18 : _GEN_369; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_371 = 5'h13 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_19 : _GEN_370; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_372 = 5'h14 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_20 : _GEN_371; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_373 = 5'h15 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_21 : _GEN_372; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_374 = 5'h16 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_22 : _GEN_373; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_375 = 5'h17 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_23 : _GEN_374; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_376 = 5'h18 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_24 : _GEN_375; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_377 = 5'h19 == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_25 : _GEN_376; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_378 = 5'h1a == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_26 : _GEN_377; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_379 = 5'h1b == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_27 : _GEN_378; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_380 = 5'h1c == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_28 : _GEN_379; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_381 = 5'h1d == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_29 : _GEN_380; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_382 = 5'h1e == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_30 : _GEN_381; // @[SIMD_ISU.scala 169:{82,82}]
  wire [4:0] _GEN_383 = 5'h1f == io_in_1_bits_ctrl_rfSrc3 ? InstBoard_io_RInstNo_31 : _GEN_382; // @[SIMD_ISU.scala 169:{82,82}]
  wire  _T_868 = _GEN_383 == io_forward_0_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_872 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_0_wb_rfDest & forwardRfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  _T_873 = _T_868 & _T_872; // @[SIMD_ISU.scala 259:140]
  wire  _T_874 = _GEN_383 == io_forward_1_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_878 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_1_wb_rfDest & forwardRfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  _T_879 = _T_874 & _T_878; // @[SIMD_ISU.scala 259:140]
  wire  _T_880 = _GEN_383 == io_forward_2_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_884 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_2_wb_rfDest & forwardRfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  _T_885 = _T_880 & _T_884; // @[SIMD_ISU.scala 259:140]
  wire  _T_886 = _GEN_383 == io_forward_3_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_890 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_3_wb_rfDest & forwardRfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  _T_891 = _T_886 & _T_890; // @[SIMD_ISU.scala 259:140]
  wire  _T_892 = _GEN_383 == io_forward_4_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_896 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_4_wb_rfDest & forwardRfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  _T_897 = _T_892 & _T_896; // @[SIMD_ISU.scala 259:140]
  wire  _T_898 = _GEN_383 == io_forward_5_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_902 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_5_wb_rfDest & forwardRfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  _T_903 = _T_898 & _T_902; // @[SIMD_ISU.scala 259:140]
  wire  _T_904 = _GEN_383 == io_forward_6_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_908 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_6_wb_rfDest & forwardRfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  _T_909 = _T_904 & _T_908; // @[SIMD_ISU.scala 259:140]
  wire  _T_910 = _GEN_383 == io_forward_7_InstNo; // @[SIMD_ISU.scala 169:82]
  wire  _T_914 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_forward_7_wb_rfDest & forwardRfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  _T_915 = _T_910 & _T_914; // @[SIMD_ISU.scala 259:140]
  wire  _T_1036 = _T_873 | _T_879 | _T_885 | _T_891 | _T_897 | _T_903 | _T_909 | _T_915; // @[SIMD_ISU.scala 261:105]
  wire  _T_964 = _GEN_383 == io_wb_InstNo_0; // @[SIMD_ISU.scala 169:82]
  wire  _T_968 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_0 & io_wb_rfWen_0; // @[SIMD_ISU.scala 166:102]
  wire  _T_969 = _T_964 & _T_968; // @[SIMD_ISU.scala 260:135]
  wire  _T_970 = _GEN_383 == io_wb_InstNo_1; // @[SIMD_ISU.scala 169:82]
  wire  _T_974 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_1 & io_wb_rfWen_1; // @[SIMD_ISU.scala 166:102]
  wire  _T_975 = _T_970 & _T_974; // @[SIMD_ISU.scala 260:135]
  wire  _T_976 = _GEN_383 == io_wb_InstNo_2; // @[SIMD_ISU.scala 169:82]
  wire  _T_980 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_2 & io_wb_rfWen_2; // @[SIMD_ISU.scala 166:102]
  wire  _T_981 = _T_976 & _T_980; // @[SIMD_ISU.scala 260:135]
  wire  _T_982 = _GEN_383 == io_wb_InstNo_3; // @[SIMD_ISU.scala 169:82]
  wire  _T_986 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_3 & io_wb_rfWen_3; // @[SIMD_ISU.scala 166:102]
  wire  _T_987 = _T_982 & _T_986; // @[SIMD_ISU.scala 260:135]
  wire  _T_988 = _GEN_383 == io_wb_InstNo_4; // @[SIMD_ISU.scala 169:82]
  wire  _T_992 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_4 & io_wb_rfWen_4; // @[SIMD_ISU.scala 166:102]
  wire  _T_993 = _T_988 & _T_992; // @[SIMD_ISU.scala 260:135]
  wire  _T_994 = _GEN_383 == io_wb_InstNo_5; // @[SIMD_ISU.scala 169:82]
  wire  _T_998 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_5 & io_wb_rfWen_5; // @[SIMD_ISU.scala 166:102]
  wire  _T_999 = _T_994 & _T_998; // @[SIMD_ISU.scala 260:135]
  wire  _T_1000 = _GEN_383 == io_wb_InstNo_6; // @[SIMD_ISU.scala 169:82]
  wire  _T_1004 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_6 & io_wb_rfWen_6; // @[SIMD_ISU.scala 166:102]
  wire  _T_1005 = _T_1000 & _T_1004; // @[SIMD_ISU.scala 260:135]
  wire  _T_1006 = _GEN_383 == io_wb_InstNo_7; // @[SIMD_ISU.scala 169:82]
  wire  _T_1010 = io_in_1_bits_ctrl_rfSrc3 != 5'h0 & io_in_1_bits_ctrl_rfSrc3 == io_wb_rfDest_7 & io_wb_rfWen_7; // @[SIMD_ISU.scala 166:102]
  wire  _T_1011 = _T_1006 & _T_1010; // @[SIMD_ISU.scala 260:135]
  wire  _T_1044 = _T_969 | _T_975 | _T_981 | _T_987 | _T_993 | _T_999 | _T_1005 | _T_1011; // @[SIMD_ISU.scala 261:135]
  wire  src3Ready_1 = ~_GEN_447 | (_T_873 | _T_879 | _T_885 | _T_891 | _T_897 | _T_903 | _T_909 | _T_915) | (_T_969 |
    _T_975 | _T_981 | _T_987 | _T_993 | _T_999 | _T_1005 | _T_1011); // @[SIMD_ISU.scala 261:109]
  wire  _T_505 = io_in_1_bits_ctrl_fuType == 4'h1 | io_in_1_bits_ctrl_fuType == 4'h8; // @[SIMD_ISU.scala 167:75]
  wire  _T_521 = io_out_0_ready & io_out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_524 = io_out_1_ready & io_out_1_valid; // @[Decoupled.scala 40:37]
  wire [24:0] _T_529 = io_in_0_bits_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_530 = {_T_529,io_in_0_bits_cf_pc}; // @[Cat.scala 30:58]
  wire [2:0] _T_538 = src1DependEX_0_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_539 = src1DependEX_0_5 ? 3'h5 : _T_538; // @[Mux.scala 47:69]
  wire [2:0] _T_540 = src1DependEX_0_4 ? 3'h4 : _T_539; // @[Mux.scala 47:69]
  wire [2:0] _T_541 = src1DependEX_0_3 ? 3'h3 : _T_540; // @[Mux.scala 47:69]
  wire [2:0] _T_542 = src1DependEX_0_2 ? 3'h2 : _T_541; // @[Mux.scala 47:69]
  wire [2:0] _T_543 = src1DependEX_0_1 ? 3'h1 : _T_542; // @[Mux.scala 47:69]
  wire [2:0] _T_544 = src1DependEX_0_0 ? 3'h0 : _T_543; // @[Mux.scala 47:69]
  wire  _T_559 = ~_T_399; // @[SIMD_ISU.scala 233:42]
  wire  _T_560 = _T_407 & ~_T_399; // @[SIMD_ISU.scala 233:39]
  wire [2:0] _T_561 = src1DependWB_0_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_562 = src1DependWB_0_5 ? 3'h5 : _T_561; // @[Mux.scala 47:69]
  wire [2:0] _T_563 = src1DependWB_0_4 ? 3'h4 : _T_562; // @[Mux.scala 47:69]
  wire [2:0] _T_564 = src1DependWB_0_3 ? 3'h3 : _T_563; // @[Mux.scala 47:69]
  wire [2:0] _T_565 = src1DependWB_0_2 ? 3'h2 : _T_564; // @[Mux.scala 47:69]
  wire [2:0] _T_566 = src1DependWB_0_1 ? 3'h1 : _T_565; // @[Mux.scala 47:69]
  wire [2:0] _T_567 = src1DependWB_0_0 ? 3'h0 : _T_566; // @[Mux.scala 47:69]
  wire  _T_586 = ~io_in_0_bits_ctrl_src1Type & _T_559 & ~_T_407; // @[SIMD_ISU.scala 234:88]
  wire [63:0] _T_587 = io_in_0_bits_ctrl_src1Type ? _T_530 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_257 = 3'h1 == _T_544 ? io_forward_1_wb_rfData : io_forward_0_wb_rfData; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_258 = 3'h2 == _T_544 ? io_forward_2_wb_rfData : _GEN_257; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_259 = 3'h3 == _T_544 ? io_forward_3_wb_rfData : _GEN_258; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_260 = 3'h4 == _T_544 ? io_forward_4_wb_rfData : _GEN_259; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_261 = 3'h5 == _T_544 ? io_forward_5_wb_rfData : _GEN_260; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_262 = 3'h6 == _T_544 ? io_forward_6_wb_rfData : _GEN_261; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_263 = 3'h7 == _T_544 ? io_forward_7_wb_rfData : _GEN_262; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_588 = _T_399 ? _GEN_263 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_265 = 3'h1 == _T_567 ? io_wb_WriteData_1 : io_wb_WriteData_0; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_266 = 3'h2 == _T_567 ? io_wb_WriteData_2 : _GEN_265; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_267 = 3'h3 == _T_567 ? io_wb_WriteData_3 : _GEN_266; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_268 = 3'h4 == _T_567 ? io_wb_WriteData_4 : _GEN_267; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_269 = 3'h5 == _T_567 ? io_wb_WriteData_5 : _GEN_268; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_270 = 3'h6 == _T_567 ? io_wb_WriteData_6 : _GEN_269; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_271 = 3'h7 == _T_567 ? io_wb_WriteData_7 : _GEN_270; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_589 = _T_560 ? _GEN_271 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_590 = _T_586 ? io_wb_ReadData1_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_591 = _T_587 | _T_588; // @[Mux.scala 27:72]
  wire [63:0] _T_592 = _T_591 | _T_589; // @[Mux.scala 27:72]
  wire [24:0] _T_597 = io_in_1_bits_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_598 = {_T_597,io_in_1_bits_cf_pc}; // @[Cat.scala 30:58]
  wire [2:0] _T_606 = src1DependEX_1_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_607 = src1DependEX_1_5 ? 3'h5 : _T_606; // @[Mux.scala 47:69]
  wire [2:0] _T_608 = src1DependEX_1_4 ? 3'h4 : _T_607; // @[Mux.scala 47:69]
  wire [2:0] _T_609 = src1DependEX_1_3 ? 3'h3 : _T_608; // @[Mux.scala 47:69]
  wire [2:0] _T_610 = src1DependEX_1_2 ? 3'h2 : _T_609; // @[Mux.scala 47:69]
  wire [2:0] _T_611 = src1DependEX_1_1 ? 3'h1 : _T_610; // @[Mux.scala 47:69]
  wire [2:0] _T_612 = src1DependEX_1_0 ? 3'h0 : _T_611; // @[Mux.scala 47:69]
  wire  _T_627 = ~_T_416; // @[SIMD_ISU.scala 233:42]
  wire  _T_628 = _T_424 & ~_T_416; // @[SIMD_ISU.scala 233:39]
  wire [2:0] _T_629 = src1DependWB_1_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_630 = src1DependWB_1_5 ? 3'h5 : _T_629; // @[Mux.scala 47:69]
  wire [2:0] _T_631 = src1DependWB_1_4 ? 3'h4 : _T_630; // @[Mux.scala 47:69]
  wire [2:0] _T_632 = src1DependWB_1_3 ? 3'h3 : _T_631; // @[Mux.scala 47:69]
  wire [2:0] _T_633 = src1DependWB_1_2 ? 3'h2 : _T_632; // @[Mux.scala 47:69]
  wire [2:0] _T_634 = src1DependWB_1_1 ? 3'h1 : _T_633; // @[Mux.scala 47:69]
  wire [2:0] _T_635 = src1DependWB_1_0 ? 3'h0 : _T_634; // @[Mux.scala 47:69]
  wire  _T_654 = ~io_in_1_bits_ctrl_src1Type & _T_627 & ~_T_424; // @[SIMD_ISU.scala 234:88]
  wire [63:0] _T_655 = io_in_1_bits_ctrl_src1Type ? _T_598 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_273 = 3'h1 == _T_612 ? io_forward_1_wb_rfData : io_forward_0_wb_rfData; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_274 = 3'h2 == _T_612 ? io_forward_2_wb_rfData : _GEN_273; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_275 = 3'h3 == _T_612 ? io_forward_3_wb_rfData : _GEN_274; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_276 = 3'h4 == _T_612 ? io_forward_4_wb_rfData : _GEN_275; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_277 = 3'h5 == _T_612 ? io_forward_5_wb_rfData : _GEN_276; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_278 = 3'h6 == _T_612 ? io_forward_6_wb_rfData : _GEN_277; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_279 = 3'h7 == _T_612 ? io_forward_7_wb_rfData : _GEN_278; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_656 = _T_416 ? _GEN_279 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_281 = 3'h1 == _T_635 ? io_wb_WriteData_1 : io_wb_WriteData_0; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_282 = 3'h2 == _T_635 ? io_wb_WriteData_2 : _GEN_281; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_283 = 3'h3 == _T_635 ? io_wb_WriteData_3 : _GEN_282; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_284 = 3'h4 == _T_635 ? io_wb_WriteData_4 : _GEN_283; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_285 = 3'h5 == _T_635 ? io_wb_WriteData_5 : _GEN_284; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_286 = 3'h6 == _T_635 ? io_wb_WriteData_6 : _GEN_285; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_287 = 3'h7 == _T_635 ? io_wb_WriteData_7 : _GEN_286; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_657 = _T_628 ? _GEN_287 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_658 = _T_654 ? io_wb_ReadData1_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_659 = _T_655 | _T_656; // @[Mux.scala 27:72]
  wire [63:0] _T_660 = _T_659 | _T_657; // @[Mux.scala 27:72]
  wire [2:0] _T_670 = src2DependEX_0_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_671 = src2DependEX_0_5 ? 3'h5 : _T_670; // @[Mux.scala 47:69]
  wire [2:0] _T_672 = src2DependEX_0_4 ? 3'h4 : _T_671; // @[Mux.scala 47:69]
  wire [2:0] _T_673 = src2DependEX_0_3 ? 3'h3 : _T_672; // @[Mux.scala 47:69]
  wire [2:0] _T_674 = src2DependEX_0_2 ? 3'h2 : _T_673; // @[Mux.scala 47:69]
  wire [2:0] _T_675 = src2DependEX_0_1 ? 3'h1 : _T_674; // @[Mux.scala 47:69]
  wire [2:0] _T_676 = src2DependEX_0_0 ? 3'h0 : _T_675; // @[Mux.scala 47:69]
  wire  _T_691 = ~_T_433; // @[SIMD_ISU.scala 241:42]
  wire  _T_692 = _T_441 & ~_T_433; // @[SIMD_ISU.scala 241:39]
  wire [2:0] _T_693 = src2DependWB_0_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_694 = src2DependWB_0_5 ? 3'h5 : _T_693; // @[Mux.scala 47:69]
  wire [2:0] _T_695 = src2DependWB_0_4 ? 3'h4 : _T_694; // @[Mux.scala 47:69]
  wire [2:0] _T_696 = src2DependWB_0_3 ? 3'h3 : _T_695; // @[Mux.scala 47:69]
  wire [2:0] _T_697 = src2DependWB_0_2 ? 3'h2 : _T_696; // @[Mux.scala 47:69]
  wire [2:0] _T_698 = src2DependWB_0_1 ? 3'h1 : _T_697; // @[Mux.scala 47:69]
  wire [2:0] _T_699 = src2DependWB_0_0 ? 3'h0 : _T_698; // @[Mux.scala 47:69]
  wire  _T_718 = ~io_in_0_bits_ctrl_src2Type & _T_691 & ~_T_441; // @[SIMD_ISU.scala 242:89]
  wire [63:0] _T_719 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_289 = 3'h1 == _T_676 ? io_forward_1_wb_rfData : io_forward_0_wb_rfData; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_290 = 3'h2 == _T_676 ? io_forward_2_wb_rfData : _GEN_289; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_291 = 3'h3 == _T_676 ? io_forward_3_wb_rfData : _GEN_290; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_292 = 3'h4 == _T_676 ? io_forward_4_wb_rfData : _GEN_291; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_293 = 3'h5 == _T_676 ? io_forward_5_wb_rfData : _GEN_292; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_294 = 3'h6 == _T_676 ? io_forward_6_wb_rfData : _GEN_293; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_295 = 3'h7 == _T_676 ? io_forward_7_wb_rfData : _GEN_294; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_720 = _T_433 ? _GEN_295 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_297 = 3'h1 == _T_699 ? io_wb_WriteData_1 : io_wb_WriteData_0; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_298 = 3'h2 == _T_699 ? io_wb_WriteData_2 : _GEN_297; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_299 = 3'h3 == _T_699 ? io_wb_WriteData_3 : _GEN_298; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_300 = 3'h4 == _T_699 ? io_wb_WriteData_4 : _GEN_299; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_301 = 3'h5 == _T_699 ? io_wb_WriteData_5 : _GEN_300; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_302 = 3'h6 == _T_699 ? io_wb_WriteData_6 : _GEN_301; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_303 = 3'h7 == _T_699 ? io_wb_WriteData_7 : _GEN_302; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_721 = _T_692 ? _GEN_303 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_722 = _T_718 ? io_wb_ReadData2_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_723 = _T_719 | _T_720; // @[Mux.scala 27:72]
  wire [63:0] _T_724 = _T_723 | _T_721; // @[Mux.scala 27:72]
  wire [2:0] _T_734 = src2DependEX_1_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_735 = src2DependEX_1_5 ? 3'h5 : _T_734; // @[Mux.scala 47:69]
  wire [2:0] _T_736 = src2DependEX_1_4 ? 3'h4 : _T_735; // @[Mux.scala 47:69]
  wire [2:0] _T_737 = src2DependEX_1_3 ? 3'h3 : _T_736; // @[Mux.scala 47:69]
  wire [2:0] _T_738 = src2DependEX_1_2 ? 3'h2 : _T_737; // @[Mux.scala 47:69]
  wire [2:0] _T_739 = src2DependEX_1_1 ? 3'h1 : _T_738; // @[Mux.scala 47:69]
  wire [2:0] _T_740 = src2DependEX_1_0 ? 3'h0 : _T_739; // @[Mux.scala 47:69]
  wire  _T_755 = ~_T_450; // @[SIMD_ISU.scala 241:42]
  wire  _T_756 = _T_458 & ~_T_450; // @[SIMD_ISU.scala 241:39]
  wire [2:0] _T_757 = src2DependWB_1_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_758 = src2DependWB_1_5 ? 3'h5 : _T_757; // @[Mux.scala 47:69]
  wire [2:0] _T_759 = src2DependWB_1_4 ? 3'h4 : _T_758; // @[Mux.scala 47:69]
  wire [2:0] _T_760 = src2DependWB_1_3 ? 3'h3 : _T_759; // @[Mux.scala 47:69]
  wire [2:0] _T_761 = src2DependWB_1_2 ? 3'h2 : _T_760; // @[Mux.scala 47:69]
  wire [2:0] _T_762 = src2DependWB_1_1 ? 3'h1 : _T_761; // @[Mux.scala 47:69]
  wire [2:0] _T_763 = src2DependWB_1_0 ? 3'h0 : _T_762; // @[Mux.scala 47:69]
  wire  _T_782 = ~io_in_1_bits_ctrl_src2Type & _T_755 & ~_T_458; // @[SIMD_ISU.scala 242:89]
  wire [63:0] _T_783 = io_in_1_bits_ctrl_src2Type ? io_in_1_bits_data_imm : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_305 = 3'h1 == _T_740 ? io_forward_1_wb_rfData : io_forward_0_wb_rfData; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_306 = 3'h2 == _T_740 ? io_forward_2_wb_rfData : _GEN_305; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_307 = 3'h3 == _T_740 ? io_forward_3_wb_rfData : _GEN_306; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_308 = 3'h4 == _T_740 ? io_forward_4_wb_rfData : _GEN_307; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_309 = 3'h5 == _T_740 ? io_forward_5_wb_rfData : _GEN_308; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_310 = 3'h6 == _T_740 ? io_forward_6_wb_rfData : _GEN_309; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_311 = 3'h7 == _T_740 ? io_forward_7_wb_rfData : _GEN_310; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_784 = _T_450 ? _GEN_311 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_313 = 3'h1 == _T_763 ? io_wb_WriteData_1 : io_wb_WriteData_0; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_314 = 3'h2 == _T_763 ? io_wb_WriteData_2 : _GEN_313; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_315 = 3'h3 == _T_763 ? io_wb_WriteData_3 : _GEN_314; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_316 = 3'h4 == _T_763 ? io_wb_WriteData_4 : _GEN_315; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_317 = 3'h5 == _T_763 ? io_wb_WriteData_5 : _GEN_316; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_318 = 3'h6 == _T_763 ? io_wb_WriteData_6 : _GEN_317; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_319 = 3'h7 == _T_763 ? io_wb_WriteData_7 : _GEN_318; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_785 = _T_756 ? _GEN_319 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_786 = _T_782 ? io_wb_ReadData2_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_787 = _T_783 | _T_784; // @[Mux.scala 27:72]
  wire [63:0] _T_788 = _T_787 | _T_785; // @[Mux.scala 27:72]
  wire [2:0] _T_1053 = _T_861 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_1054 = _T_855 ? 3'h5 : _T_1053; // @[Mux.scala 47:69]
  wire [2:0] _T_1055 = _T_849 ? 3'h4 : _T_1054; // @[Mux.scala 47:69]
  wire [2:0] _T_1056 = _T_843 ? 3'h3 : _T_1055; // @[Mux.scala 47:69]
  wire [2:0] _T_1057 = _T_837 ? 3'h2 : _T_1056; // @[Mux.scala 47:69]
  wire [2:0] _T_1058 = _T_831 ? 3'h1 : _T_1057; // @[Mux.scala 47:69]
  wire [2:0] _T_1059 = _T_825 ? 3'h0 : _T_1058; // @[Mux.scala 47:69]
  wire  _T_1074 = ~_T_1019; // @[SIMD_ISU.scala 265:42]
  wire  _T_1075 = _T_1027 & ~_T_1019; // @[SIMD_ISU.scala 265:39]
  wire [2:0] _T_1076 = _T_957 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_1077 = _T_951 ? 3'h5 : _T_1076; // @[Mux.scala 47:69]
  wire [2:0] _T_1078 = _T_945 ? 3'h4 : _T_1077; // @[Mux.scala 47:69]
  wire [2:0] _T_1079 = _T_939 ? 3'h3 : _T_1078; // @[Mux.scala 47:69]
  wire [2:0] _T_1080 = _T_933 ? 3'h2 : _T_1079; // @[Mux.scala 47:69]
  wire [2:0] _T_1081 = _T_927 ? 3'h1 : _T_1080; // @[Mux.scala 47:69]
  wire [2:0] _T_1082 = _T_921 ? 3'h0 : _T_1081; // @[Mux.scala 47:69]
  wire  _T_1099 = _T_1074 & ~_T_1027; // @[SIMD_ISU.scala 266:40]
  wire [63:0] _GEN_449 = 3'h1 == _T_1059 ? io_forward_1_wb_rfData : io_forward_0_wb_rfData; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_450 = 3'h2 == _T_1059 ? io_forward_2_wb_rfData : _GEN_449; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_451 = 3'h3 == _T_1059 ? io_forward_3_wb_rfData : _GEN_450; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_452 = 3'h4 == _T_1059 ? io_forward_4_wb_rfData : _GEN_451; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_453 = 3'h5 == _T_1059 ? io_forward_5_wb_rfData : _GEN_452; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_454 = 3'h6 == _T_1059 ? io_forward_6_wb_rfData : _GEN_453; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_455 = 3'h7 == _T_1059 ? io_forward_7_wb_rfData : _GEN_454; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_1100 = _T_1019 ? _GEN_455 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_457 = 3'h1 == _T_1082 ? io_wb_WriteData_1 : io_wb_WriteData_0; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_458 = 3'h2 == _T_1082 ? io_wb_WriteData_2 : _GEN_457; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_459 = 3'h3 == _T_1082 ? io_wb_WriteData_3 : _GEN_458; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_460 = 3'h4 == _T_1082 ? io_wb_WriteData_4 : _GEN_459; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_461 = 3'h5 == _T_1082 ? io_wb_WriteData_5 : _GEN_460; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_462 = 3'h6 == _T_1082 ? io_wb_WriteData_6 : _GEN_461; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_463 = 3'h7 == _T_1082 ? io_wb_WriteData_7 : _GEN_462; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_1101 = _T_1075 ? _GEN_463 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1102 = _T_1099 ? io_wb_ReadData3_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1103 = _T_1100 | _T_1101; // @[Mux.scala 27:72]
  wire [2:0] _T_1112 = _T_909 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_1113 = _T_903 ? 3'h5 : _T_1112; // @[Mux.scala 47:69]
  wire [2:0] _T_1114 = _T_897 ? 3'h4 : _T_1113; // @[Mux.scala 47:69]
  wire [2:0] _T_1115 = _T_891 ? 3'h3 : _T_1114; // @[Mux.scala 47:69]
  wire [2:0] _T_1116 = _T_885 ? 3'h2 : _T_1115; // @[Mux.scala 47:69]
  wire [2:0] _T_1117 = _T_879 ? 3'h1 : _T_1116; // @[Mux.scala 47:69]
  wire [2:0] _T_1118 = _T_873 ? 3'h0 : _T_1117; // @[Mux.scala 47:69]
  wire  _T_1133 = ~_T_1036; // @[SIMD_ISU.scala 265:42]
  wire  _T_1134 = _T_1044 & ~_T_1036; // @[SIMD_ISU.scala 265:39]
  wire [2:0] _T_1135 = _T_1005 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_1136 = _T_999 ? 3'h5 : _T_1135; // @[Mux.scala 47:69]
  wire [2:0] _T_1137 = _T_993 ? 3'h4 : _T_1136; // @[Mux.scala 47:69]
  wire [2:0] _T_1138 = _T_987 ? 3'h3 : _T_1137; // @[Mux.scala 47:69]
  wire [2:0] _T_1139 = _T_981 ? 3'h2 : _T_1138; // @[Mux.scala 47:69]
  wire [2:0] _T_1140 = _T_975 ? 3'h1 : _T_1139; // @[Mux.scala 47:69]
  wire [2:0] _T_1141 = _T_969 ? 3'h0 : _T_1140; // @[Mux.scala 47:69]
  wire  _T_1158 = _T_1133 & ~_T_1044; // @[SIMD_ISU.scala 266:40]
  wire [63:0] _GEN_465 = 3'h1 == _T_1118 ? io_forward_1_wb_rfData : io_forward_0_wb_rfData; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_466 = 3'h2 == _T_1118 ? io_forward_2_wb_rfData : _GEN_465; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_467 = 3'h3 == _T_1118 ? io_forward_3_wb_rfData : _GEN_466; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_468 = 3'h4 == _T_1118 ? io_forward_4_wb_rfData : _GEN_467; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_469 = 3'h5 == _T_1118 ? io_forward_5_wb_rfData : _GEN_468; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_470 = 3'h6 == _T_1118 ? io_forward_6_wb_rfData : _GEN_469; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_471 = 3'h7 == _T_1118 ? io_forward_7_wb_rfData : _GEN_470; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_1159 = _T_1036 ? _GEN_471 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_473 = 3'h1 == _T_1141 ? io_wb_WriteData_1 : io_wb_WriteData_0; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_474 = 3'h2 == _T_1141 ? io_wb_WriteData_2 : _GEN_473; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_475 = 3'h3 == _T_1141 ? io_wb_WriteData_3 : _GEN_474; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_476 = 3'h4 == _T_1141 ? io_wb_WriteData_4 : _GEN_475; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_477 = 3'h5 == _T_1141 ? io_wb_WriteData_5 : _GEN_476; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_478 = 3'h6 == _T_1141 ? io_wb_WriteData_6 : _GEN_477; // @[Mux.scala 27:{72,72}]
  wire [63:0] _GEN_479 = 3'h7 == _T_1141 ? io_wb_WriteData_7 : _GEN_478; // @[Mux.scala 27:{72,72}]
  wire [63:0] _T_1160 = _T_1134 ? _GEN_479 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1161 = _T_1158 ? io_wb_ReadData3_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1162 = _T_1159 | _T_1160; // @[Mux.scala 27:72]
  wire [1:0] _T_1166 = _T_521 + _T_524; // @[SIMD_ISU.scala 272:61]
  wire [5:0] _T_1167 = {{1'd0}, q_io_HeadPtr}; // @[SIMD_ISU.scala 276:42]
  wire  _T_1168 = _T_1167 >= 6'h20; // @[SIMD_ISU.scala 277:43]
  wire [5:0] _T_1170 = _T_1167 - 6'h20; // @[SIMD_ISU.scala 278:65]
  wire [5:0] _T_1171 = _T_1168 ? _T_1170 : _T_1167; // @[SIMD_ISU.scala 278:37]
  wire [5:0] _T_1174 = q_io_HeadPtr + 5'h1; // @[SIMD_ISU.scala 276:42]
  wire  _T_1175 = _T_1174 >= 6'h20; // @[SIMD_ISU.scala 277:43]
  wire [5:0] _T_1177 = _T_1174 - 6'h20; // @[SIMD_ISU.scala 278:65]
  wire [5:0] _T_1178 = _T_1175 ? _T_1177 : _T_1174; // @[SIMD_ISU.scala 278:37]
  wire  _T_1193 = 5'h1 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1197 = 5'h1 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1202 = 5'h2 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1206 = 5'h2 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1211 = 5'h3 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1215 = 5'h3 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1220 = 5'h4 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1224 = 5'h4 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1229 = 5'h5 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1233 = 5'h5 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1238 = 5'h6 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1242 = 5'h6 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1247 = 5'h7 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1251 = 5'h7 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1256 = 5'h8 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1260 = 5'h8 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1265 = 5'h9 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1269 = 5'h9 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1274 = 5'ha == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1278 = 5'ha == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1283 = 5'hb == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1287 = 5'hb == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1292 = 5'hc == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1296 = 5'hc == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1301 = 5'hd == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1305 = 5'hd == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1310 = 5'he == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1314 = 5'he == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1319 = 5'hf == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1323 = 5'hf == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1328 = 5'h10 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1332 = 5'h10 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1337 = 5'h11 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1341 = 5'h11 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1346 = 5'h12 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1350 = 5'h12 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1355 = 5'h13 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1359 = 5'h13 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1364 = 5'h14 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1368 = 5'h14 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1373 = 5'h15 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1377 = 5'h15 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1382 = 5'h16 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1386 = 5'h16 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1391 = 5'h17 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1395 = 5'h17 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1400 = 5'h18 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1404 = 5'h18 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1409 = 5'h19 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1413 = 5'h19 == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1418 = 5'h1a == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1422 = 5'h1a == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1427 = 5'h1b == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1431 = 5'h1b == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1436 = 5'h1c == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1440 = 5'h1c == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1445 = 5'h1d == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1449 = 5'h1d == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1454 = 5'h1e == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1458 = 5'h1e == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1463 = 5'h1f == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire  _T_1467 = 5'h1f == io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:132]
  wire [4:0] _GEN_482 = _T_1193 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_484 = _T_1202 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_486 = _T_1211 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_488 = _T_1220 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_490 = _T_1229 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_492 = _T_1238 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_494 = _T_1247 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_496 = _T_1256 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_498 = _T_1265 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_500 = _T_1274 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_502 = _T_1283 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_504 = _T_1292 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_506 = _T_1301 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_508 = _T_1310 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_510 = _T_1319 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_512 = _T_1328 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_514 = _T_1337 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_516 = _T_1346 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_518 = _T_1355 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_520 = _T_1364 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_522 = _T_1373 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_524 = _T_1382 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_526 = _T_1391 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_528 = _T_1400 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_530 = _T_1409 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_532 = _T_1418 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_534 = _T_1427 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_536 = _T_1436 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_538 = _T_1445 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_540 = _T_1454 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire [4:0] _GEN_542 = _T_1463 ? io_out_0_bits_InstNo : 5'h0; // @[SIMD_ISU.scala 287:116 285:69 288:73]
  wire  _T_1791 = io_wb_rfWen_6 & 5'h1 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_1; // @[SIMD_ISU.scala 291:140]
  wire  _T_1801 = io_wb_rfWen_0 & 5'h1 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_1 | io_wb_rfWen_1 & 5'h1
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_1 | io_wb_rfWen_2 & 5'h1 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_1 | io_wb_rfWen_3 & 5'h1 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_1 | io_wb_rfWen_4 & 5'h1 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_1 |
    io_wb_rfWen_5 & 5'h1 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_1 | _T_1791; // @[SIMD_ISU.scala 291:197]
  wire  _T_1830 = io_wb_rfWen_6 & 5'h2 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_2; // @[SIMD_ISU.scala 291:140]
  wire  _T_1840 = io_wb_rfWen_0 & 5'h2 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_2 | io_wb_rfWen_1 & 5'h2
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_2 | io_wb_rfWen_2 & 5'h2 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_2 | io_wb_rfWen_3 & 5'h2 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_2 | io_wb_rfWen_4 & 5'h2 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_2 |
    io_wb_rfWen_5 & 5'h2 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_2 | _T_1830; // @[SIMD_ISU.scala 291:197]
  wire  _T_1869 = io_wb_rfWen_6 & 5'h3 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_3; // @[SIMD_ISU.scala 291:140]
  wire  _T_1879 = io_wb_rfWen_0 & 5'h3 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_3 | io_wb_rfWen_1 & 5'h3
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_3 | io_wb_rfWen_2 & 5'h3 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_3 | io_wb_rfWen_3 & 5'h3 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_3 | io_wb_rfWen_4 & 5'h3 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_3 |
    io_wb_rfWen_5 & 5'h3 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_3 | _T_1869; // @[SIMD_ISU.scala 291:197]
  wire  _T_1908 = io_wb_rfWen_6 & 5'h4 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_4; // @[SIMD_ISU.scala 291:140]
  wire  _T_1918 = io_wb_rfWen_0 & 5'h4 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_4 | io_wb_rfWen_1 & 5'h4
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_4 | io_wb_rfWen_2 & 5'h4 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_4 | io_wb_rfWen_3 & 5'h4 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_4 | io_wb_rfWen_4 & 5'h4 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_4 |
    io_wb_rfWen_5 & 5'h4 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_4 | _T_1908; // @[SIMD_ISU.scala 291:197]
  wire  _T_1947 = io_wb_rfWen_6 & 5'h5 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_5; // @[SIMD_ISU.scala 291:140]
  wire  _T_1957 = io_wb_rfWen_0 & 5'h5 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_5 | io_wb_rfWen_1 & 5'h5
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_5 | io_wb_rfWen_2 & 5'h5 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_5 | io_wb_rfWen_3 & 5'h5 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_5 | io_wb_rfWen_4 & 5'h5 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_5 |
    io_wb_rfWen_5 & 5'h5 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_5 | _T_1947; // @[SIMD_ISU.scala 291:197]
  wire  _T_1986 = io_wb_rfWen_6 & 5'h6 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_6; // @[SIMD_ISU.scala 291:140]
  wire  _T_1996 = io_wb_rfWen_0 & 5'h6 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_6 | io_wb_rfWen_1 & 5'h6
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_6 | io_wb_rfWen_2 & 5'h6 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_6 | io_wb_rfWen_3 & 5'h6 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_6 | io_wb_rfWen_4 & 5'h6 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_6 |
    io_wb_rfWen_5 & 5'h6 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_6 | _T_1986; // @[SIMD_ISU.scala 291:197]
  wire  _T_2025 = io_wb_rfWen_6 & 5'h7 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_7; // @[SIMD_ISU.scala 291:140]
  wire  _T_2035 = io_wb_rfWen_0 & 5'h7 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_7 | io_wb_rfWen_1 & 5'h7
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_7 | io_wb_rfWen_2 & 5'h7 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_7 | io_wb_rfWen_3 & 5'h7 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_7 | io_wb_rfWen_4 & 5'h7 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_7 |
    io_wb_rfWen_5 & 5'h7 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_7 | _T_2025; // @[SIMD_ISU.scala 291:197]
  wire  _T_2064 = io_wb_rfWen_6 & 5'h8 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_8; // @[SIMD_ISU.scala 291:140]
  wire  _T_2074 = io_wb_rfWen_0 & 5'h8 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_8 | io_wb_rfWen_1 & 5'h8
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_8 | io_wb_rfWen_2 & 5'h8 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_8 | io_wb_rfWen_3 & 5'h8 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_8 | io_wb_rfWen_4 & 5'h8 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_8 |
    io_wb_rfWen_5 & 5'h8 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_8 | _T_2064; // @[SIMD_ISU.scala 291:197]
  wire  _T_2103 = io_wb_rfWen_6 & 5'h9 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_9; // @[SIMD_ISU.scala 291:140]
  wire  _T_2113 = io_wb_rfWen_0 & 5'h9 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_9 | io_wb_rfWen_1 & 5'h9
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_9 | io_wb_rfWen_2 & 5'h9 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_9 | io_wb_rfWen_3 & 5'h9 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_9 | io_wb_rfWen_4 & 5'h9 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_9 |
    io_wb_rfWen_5 & 5'h9 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_9 | _T_2103; // @[SIMD_ISU.scala 291:197]
  wire  _T_2142 = io_wb_rfWen_6 & 5'ha == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_10; // @[SIMD_ISU.scala 291:140]
  wire  _T_2152 = io_wb_rfWen_0 & 5'ha == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_10 | io_wb_rfWen_1 & 5'ha
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_10 | io_wb_rfWen_2 & 5'ha == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_10 | io_wb_rfWen_3 & 5'ha == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_10 | io_wb_rfWen_4 & 5'ha == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_10 |
    io_wb_rfWen_5 & 5'ha == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_10 | _T_2142; // @[SIMD_ISU.scala 291:197]
  wire  _T_2181 = io_wb_rfWen_6 & 5'hb == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_11; // @[SIMD_ISU.scala 291:140]
  wire  _T_2191 = io_wb_rfWen_0 & 5'hb == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_11 | io_wb_rfWen_1 & 5'hb
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_11 | io_wb_rfWen_2 & 5'hb == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_11 | io_wb_rfWen_3 & 5'hb == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_11 | io_wb_rfWen_4 & 5'hb == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_11 |
    io_wb_rfWen_5 & 5'hb == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_11 | _T_2181; // @[SIMD_ISU.scala 291:197]
  wire  _T_2220 = io_wb_rfWen_6 & 5'hc == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_12; // @[SIMD_ISU.scala 291:140]
  wire  _T_2230 = io_wb_rfWen_0 & 5'hc == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_12 | io_wb_rfWen_1 & 5'hc
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_12 | io_wb_rfWen_2 & 5'hc == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_12 | io_wb_rfWen_3 & 5'hc == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_12 | io_wb_rfWen_4 & 5'hc == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_12 |
    io_wb_rfWen_5 & 5'hc == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_12 | _T_2220; // @[SIMD_ISU.scala 291:197]
  wire  _T_2259 = io_wb_rfWen_6 & 5'hd == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_13; // @[SIMD_ISU.scala 291:140]
  wire  _T_2269 = io_wb_rfWen_0 & 5'hd == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_13 | io_wb_rfWen_1 & 5'hd
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_13 | io_wb_rfWen_2 & 5'hd == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_13 | io_wb_rfWen_3 & 5'hd == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_13 | io_wb_rfWen_4 & 5'hd == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_13 |
    io_wb_rfWen_5 & 5'hd == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_13 | _T_2259; // @[SIMD_ISU.scala 291:197]
  wire  _T_2298 = io_wb_rfWen_6 & 5'he == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_14; // @[SIMD_ISU.scala 291:140]
  wire  _T_2308 = io_wb_rfWen_0 & 5'he == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_14 | io_wb_rfWen_1 & 5'he
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_14 | io_wb_rfWen_2 & 5'he == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_14 | io_wb_rfWen_3 & 5'he == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_14 | io_wb_rfWen_4 & 5'he == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_14 |
    io_wb_rfWen_5 & 5'he == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_14 | _T_2298; // @[SIMD_ISU.scala 291:197]
  wire  _T_2337 = io_wb_rfWen_6 & 5'hf == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_15; // @[SIMD_ISU.scala 291:140]
  wire  _T_2347 = io_wb_rfWen_0 & 5'hf == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_15 | io_wb_rfWen_1 & 5'hf
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_15 | io_wb_rfWen_2 & 5'hf == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_15 | io_wb_rfWen_3 & 5'hf == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_15 | io_wb_rfWen_4 & 5'hf == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_15 |
    io_wb_rfWen_5 & 5'hf == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_15 | _T_2337; // @[SIMD_ISU.scala 291:197]
  wire  _T_2376 = io_wb_rfWen_6 & 5'h10 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_16; // @[SIMD_ISU.scala 291:140]
  wire  _T_2386 = io_wb_rfWen_0 & 5'h10 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_16 | io_wb_rfWen_1 & 5'h10
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_16 | io_wb_rfWen_2 & 5'h10 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_16 | io_wb_rfWen_3 & 5'h10 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_16 | io_wb_rfWen_4 & 5'h10 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_16 |
    io_wb_rfWen_5 & 5'h10 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_16 | _T_2376; // @[SIMD_ISU.scala 291:197]
  wire  _T_2415 = io_wb_rfWen_6 & 5'h11 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_17; // @[SIMD_ISU.scala 291:140]
  wire  _T_2425 = io_wb_rfWen_0 & 5'h11 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_17 | io_wb_rfWen_1 & 5'h11
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_17 | io_wb_rfWen_2 & 5'h11 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_17 | io_wb_rfWen_3 & 5'h11 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_17 | io_wb_rfWen_4 & 5'h11 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_17 |
    io_wb_rfWen_5 & 5'h11 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_17 | _T_2415; // @[SIMD_ISU.scala 291:197]
  wire  _T_2454 = io_wb_rfWen_6 & 5'h12 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_18; // @[SIMD_ISU.scala 291:140]
  wire  _T_2464 = io_wb_rfWen_0 & 5'h12 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_18 | io_wb_rfWen_1 & 5'h12
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_18 | io_wb_rfWen_2 & 5'h12 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_18 | io_wb_rfWen_3 & 5'h12 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_18 | io_wb_rfWen_4 & 5'h12 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_18 |
    io_wb_rfWen_5 & 5'h12 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_18 | _T_2454; // @[SIMD_ISU.scala 291:197]
  wire  _T_2493 = io_wb_rfWen_6 & 5'h13 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_19; // @[SIMD_ISU.scala 291:140]
  wire  _T_2503 = io_wb_rfWen_0 & 5'h13 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_19 | io_wb_rfWen_1 & 5'h13
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_19 | io_wb_rfWen_2 & 5'h13 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_19 | io_wb_rfWen_3 & 5'h13 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_19 | io_wb_rfWen_4 & 5'h13 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_19 |
    io_wb_rfWen_5 & 5'h13 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_19 | _T_2493; // @[SIMD_ISU.scala 291:197]
  wire  _T_2532 = io_wb_rfWen_6 & 5'h14 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_20; // @[SIMD_ISU.scala 291:140]
  wire  _T_2542 = io_wb_rfWen_0 & 5'h14 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_20 | io_wb_rfWen_1 & 5'h14
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_20 | io_wb_rfWen_2 & 5'h14 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_20 | io_wb_rfWen_3 & 5'h14 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_20 | io_wb_rfWen_4 & 5'h14 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_20 |
    io_wb_rfWen_5 & 5'h14 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_20 | _T_2532; // @[SIMD_ISU.scala 291:197]
  wire  _T_2571 = io_wb_rfWen_6 & 5'h15 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_21; // @[SIMD_ISU.scala 291:140]
  wire  _T_2581 = io_wb_rfWen_0 & 5'h15 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_21 | io_wb_rfWen_1 & 5'h15
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_21 | io_wb_rfWen_2 & 5'h15 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_21 | io_wb_rfWen_3 & 5'h15 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_21 | io_wb_rfWen_4 & 5'h15 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_21 |
    io_wb_rfWen_5 & 5'h15 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_21 | _T_2571; // @[SIMD_ISU.scala 291:197]
  wire  _T_2610 = io_wb_rfWen_6 & 5'h16 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_22; // @[SIMD_ISU.scala 291:140]
  wire  _T_2620 = io_wb_rfWen_0 & 5'h16 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_22 | io_wb_rfWen_1 & 5'h16
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_22 | io_wb_rfWen_2 & 5'h16 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_22 | io_wb_rfWen_3 & 5'h16 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_22 | io_wb_rfWen_4 & 5'h16 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_22 |
    io_wb_rfWen_5 & 5'h16 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_22 | _T_2610; // @[SIMD_ISU.scala 291:197]
  wire  _T_2649 = io_wb_rfWen_6 & 5'h17 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_23; // @[SIMD_ISU.scala 291:140]
  wire  _T_2659 = io_wb_rfWen_0 & 5'h17 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_23 | io_wb_rfWen_1 & 5'h17
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_23 | io_wb_rfWen_2 & 5'h17 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_23 | io_wb_rfWen_3 & 5'h17 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_23 | io_wb_rfWen_4 & 5'h17 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_23 |
    io_wb_rfWen_5 & 5'h17 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_23 | _T_2649; // @[SIMD_ISU.scala 291:197]
  wire  _T_2688 = io_wb_rfWen_6 & 5'h18 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_24; // @[SIMD_ISU.scala 291:140]
  wire  _T_2698 = io_wb_rfWen_0 & 5'h18 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_24 | io_wb_rfWen_1 & 5'h18
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_24 | io_wb_rfWen_2 & 5'h18 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_24 | io_wb_rfWen_3 & 5'h18 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_24 | io_wb_rfWen_4 & 5'h18 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_24 |
    io_wb_rfWen_5 & 5'h18 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_24 | _T_2688; // @[SIMD_ISU.scala 291:197]
  wire  _T_2727 = io_wb_rfWen_6 & 5'h19 == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_25; // @[SIMD_ISU.scala 291:140]
  wire  _T_2737 = io_wb_rfWen_0 & 5'h19 == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_25 | io_wb_rfWen_1 & 5'h19
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_25 | io_wb_rfWen_2 & 5'h19 == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_25 | io_wb_rfWen_3 & 5'h19 == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_25 | io_wb_rfWen_4 & 5'h19 == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_25 |
    io_wb_rfWen_5 & 5'h19 == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_25 | _T_2727; // @[SIMD_ISU.scala 291:197]
  wire  _T_2766 = io_wb_rfWen_6 & 5'h1a == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_26; // @[SIMD_ISU.scala 291:140]
  wire  _T_2776 = io_wb_rfWen_0 & 5'h1a == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_26 | io_wb_rfWen_1 & 5'h1a
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_26 | io_wb_rfWen_2 & 5'h1a == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_26 | io_wb_rfWen_3 & 5'h1a == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_26 | io_wb_rfWen_4 & 5'h1a == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_26 |
    io_wb_rfWen_5 & 5'h1a == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_26 | _T_2766; // @[SIMD_ISU.scala 291:197]
  wire  _T_2805 = io_wb_rfWen_6 & 5'h1b == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_27; // @[SIMD_ISU.scala 291:140]
  wire  _T_2815 = io_wb_rfWen_0 & 5'h1b == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_27 | io_wb_rfWen_1 & 5'h1b
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_27 | io_wb_rfWen_2 & 5'h1b == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_27 | io_wb_rfWen_3 & 5'h1b == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_27 | io_wb_rfWen_4 & 5'h1b == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_27 |
    io_wb_rfWen_5 & 5'h1b == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_27 | _T_2805; // @[SIMD_ISU.scala 291:197]
  wire  _T_2844 = io_wb_rfWen_6 & 5'h1c == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_28; // @[SIMD_ISU.scala 291:140]
  wire  _T_2854 = io_wb_rfWen_0 & 5'h1c == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_28 | io_wb_rfWen_1 & 5'h1c
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_28 | io_wb_rfWen_2 & 5'h1c == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_28 | io_wb_rfWen_3 & 5'h1c == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_28 | io_wb_rfWen_4 & 5'h1c == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_28 |
    io_wb_rfWen_5 & 5'h1c == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_28 | _T_2844; // @[SIMD_ISU.scala 291:197]
  wire  _T_2883 = io_wb_rfWen_6 & 5'h1d == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_29; // @[SIMD_ISU.scala 291:140]
  wire  _T_2893 = io_wb_rfWen_0 & 5'h1d == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_29 | io_wb_rfWen_1 & 5'h1d
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_29 | io_wb_rfWen_2 & 5'h1d == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_29 | io_wb_rfWen_3 & 5'h1d == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_29 | io_wb_rfWen_4 & 5'h1d == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_29 |
    io_wb_rfWen_5 & 5'h1d == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_29 | _T_2883; // @[SIMD_ISU.scala 291:197]
  wire  _T_2922 = io_wb_rfWen_6 & 5'h1e == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_30; // @[SIMD_ISU.scala 291:140]
  wire  _T_2932 = io_wb_rfWen_0 & 5'h1e == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_30 | io_wb_rfWen_1 & 5'h1e
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_30 | io_wb_rfWen_2 & 5'h1e == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_30 | io_wb_rfWen_3 & 5'h1e == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_30 | io_wb_rfWen_4 & 5'h1e == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_30 |
    io_wb_rfWen_5 & 5'h1e == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_30 | _T_2922; // @[SIMD_ISU.scala 291:197]
  wire  _T_2961 = io_wb_rfWen_6 & 5'h1f == io_wb_rfDest_6 & io_wb_InstNo_6 == InstBoard_io_RInstNo_31; // @[SIMD_ISU.scala 291:140]
  wire  _T_2971 = io_wb_rfWen_0 & 5'h1f == io_wb_rfDest_0 & io_wb_InstNo_0 == InstBoard_io_RInstNo_31 | io_wb_rfWen_1 & 5'h1f
     == io_wb_rfDest_1 & io_wb_InstNo_1 == InstBoard_io_RInstNo_31 | io_wb_rfWen_2 & 5'h1f == io_wb_rfDest_2 &
    io_wb_InstNo_2 == InstBoard_io_RInstNo_31 | io_wb_rfWen_3 & 5'h1f == io_wb_rfDest_3 & io_wb_InstNo_3 ==
    InstBoard_io_RInstNo_31 | io_wb_rfWen_4 & 5'h1f == io_wb_rfDest_4 & io_wb_InstNo_4 == InstBoard_io_RInstNo_31 |
    io_wb_rfWen_5 & 5'h1f == io_wb_rfDest_5 & io_wb_InstNo_5 == InstBoard_io_RInstNo_31 | _T_2961; // @[SIMD_ISU.scala 291:197]
  InstBoard InstBoard ( // @[SIMD_ISU.scala 163:27]
    .clock(InstBoard_clock),
    .reset(InstBoard_reset),
    .io_Wen_1(InstBoard_io_Wen_1),
    .io_Wen_2(InstBoard_io_Wen_2),
    .io_Wen_3(InstBoard_io_Wen_3),
    .io_Wen_4(InstBoard_io_Wen_4),
    .io_Wen_5(InstBoard_io_Wen_5),
    .io_Wen_6(InstBoard_io_Wen_6),
    .io_Wen_7(InstBoard_io_Wen_7),
    .io_Wen_8(InstBoard_io_Wen_8),
    .io_Wen_9(InstBoard_io_Wen_9),
    .io_Wen_10(InstBoard_io_Wen_10),
    .io_Wen_11(InstBoard_io_Wen_11),
    .io_Wen_12(InstBoard_io_Wen_12),
    .io_Wen_13(InstBoard_io_Wen_13),
    .io_Wen_14(InstBoard_io_Wen_14),
    .io_Wen_15(InstBoard_io_Wen_15),
    .io_Wen_16(InstBoard_io_Wen_16),
    .io_Wen_17(InstBoard_io_Wen_17),
    .io_Wen_18(InstBoard_io_Wen_18),
    .io_Wen_19(InstBoard_io_Wen_19),
    .io_Wen_20(InstBoard_io_Wen_20),
    .io_Wen_21(InstBoard_io_Wen_21),
    .io_Wen_22(InstBoard_io_Wen_22),
    .io_Wen_23(InstBoard_io_Wen_23),
    .io_Wen_24(InstBoard_io_Wen_24),
    .io_Wen_25(InstBoard_io_Wen_25),
    .io_Wen_26(InstBoard_io_Wen_26),
    .io_Wen_27(InstBoard_io_Wen_27),
    .io_Wen_28(InstBoard_io_Wen_28),
    .io_Wen_29(InstBoard_io_Wen_29),
    .io_Wen_30(InstBoard_io_Wen_30),
    .io_Wen_31(InstBoard_io_Wen_31),
    .io_clear_1(InstBoard_io_clear_1),
    .io_clear_2(InstBoard_io_clear_2),
    .io_clear_3(InstBoard_io_clear_3),
    .io_clear_4(InstBoard_io_clear_4),
    .io_clear_5(InstBoard_io_clear_5),
    .io_clear_6(InstBoard_io_clear_6),
    .io_clear_7(InstBoard_io_clear_7),
    .io_clear_8(InstBoard_io_clear_8),
    .io_clear_9(InstBoard_io_clear_9),
    .io_clear_10(InstBoard_io_clear_10),
    .io_clear_11(InstBoard_io_clear_11),
    .io_clear_12(InstBoard_io_clear_12),
    .io_clear_13(InstBoard_io_clear_13),
    .io_clear_14(InstBoard_io_clear_14),
    .io_clear_15(InstBoard_io_clear_15),
    .io_clear_16(InstBoard_io_clear_16),
    .io_clear_17(InstBoard_io_clear_17),
    .io_clear_18(InstBoard_io_clear_18),
    .io_clear_19(InstBoard_io_clear_19),
    .io_clear_20(InstBoard_io_clear_20),
    .io_clear_21(InstBoard_io_clear_21),
    .io_clear_22(InstBoard_io_clear_22),
    .io_clear_23(InstBoard_io_clear_23),
    .io_clear_24(InstBoard_io_clear_24),
    .io_clear_25(InstBoard_io_clear_25),
    .io_clear_26(InstBoard_io_clear_26),
    .io_clear_27(InstBoard_io_clear_27),
    .io_clear_28(InstBoard_io_clear_28),
    .io_clear_29(InstBoard_io_clear_29),
    .io_clear_30(InstBoard_io_clear_30),
    .io_clear_31(InstBoard_io_clear_31),
    .io_WInstNo_1(InstBoard_io_WInstNo_1),
    .io_WInstNo_2(InstBoard_io_WInstNo_2),
    .io_WInstNo_3(InstBoard_io_WInstNo_3),
    .io_WInstNo_4(InstBoard_io_WInstNo_4),
    .io_WInstNo_5(InstBoard_io_WInstNo_5),
    .io_WInstNo_6(InstBoard_io_WInstNo_6),
    .io_WInstNo_7(InstBoard_io_WInstNo_7),
    .io_WInstNo_8(InstBoard_io_WInstNo_8),
    .io_WInstNo_9(InstBoard_io_WInstNo_9),
    .io_WInstNo_10(InstBoard_io_WInstNo_10),
    .io_WInstNo_11(InstBoard_io_WInstNo_11),
    .io_WInstNo_12(InstBoard_io_WInstNo_12),
    .io_WInstNo_13(InstBoard_io_WInstNo_13),
    .io_WInstNo_14(InstBoard_io_WInstNo_14),
    .io_WInstNo_15(InstBoard_io_WInstNo_15),
    .io_WInstNo_16(InstBoard_io_WInstNo_16),
    .io_WInstNo_17(InstBoard_io_WInstNo_17),
    .io_WInstNo_18(InstBoard_io_WInstNo_18),
    .io_WInstNo_19(InstBoard_io_WInstNo_19),
    .io_WInstNo_20(InstBoard_io_WInstNo_20),
    .io_WInstNo_21(InstBoard_io_WInstNo_21),
    .io_WInstNo_22(InstBoard_io_WInstNo_22),
    .io_WInstNo_23(InstBoard_io_WInstNo_23),
    .io_WInstNo_24(InstBoard_io_WInstNo_24),
    .io_WInstNo_25(InstBoard_io_WInstNo_25),
    .io_WInstNo_26(InstBoard_io_WInstNo_26),
    .io_WInstNo_27(InstBoard_io_WInstNo_27),
    .io_WInstNo_28(InstBoard_io_WInstNo_28),
    .io_WInstNo_29(InstBoard_io_WInstNo_29),
    .io_WInstNo_30(InstBoard_io_WInstNo_30),
    .io_WInstNo_31(InstBoard_io_WInstNo_31),
    .io_valid_1(InstBoard_io_valid_1),
    .io_valid_2(InstBoard_io_valid_2),
    .io_valid_3(InstBoard_io_valid_3),
    .io_valid_4(InstBoard_io_valid_4),
    .io_valid_5(InstBoard_io_valid_5),
    .io_valid_6(InstBoard_io_valid_6),
    .io_valid_7(InstBoard_io_valid_7),
    .io_valid_8(InstBoard_io_valid_8),
    .io_valid_9(InstBoard_io_valid_9),
    .io_valid_10(InstBoard_io_valid_10),
    .io_valid_11(InstBoard_io_valid_11),
    .io_valid_12(InstBoard_io_valid_12),
    .io_valid_13(InstBoard_io_valid_13),
    .io_valid_14(InstBoard_io_valid_14),
    .io_valid_15(InstBoard_io_valid_15),
    .io_valid_16(InstBoard_io_valid_16),
    .io_valid_17(InstBoard_io_valid_17),
    .io_valid_18(InstBoard_io_valid_18),
    .io_valid_19(InstBoard_io_valid_19),
    .io_valid_20(InstBoard_io_valid_20),
    .io_valid_21(InstBoard_io_valid_21),
    .io_valid_22(InstBoard_io_valid_22),
    .io_valid_23(InstBoard_io_valid_23),
    .io_valid_24(InstBoard_io_valid_24),
    .io_valid_25(InstBoard_io_valid_25),
    .io_valid_26(InstBoard_io_valid_26),
    .io_valid_27(InstBoard_io_valid_27),
    .io_valid_28(InstBoard_io_valid_28),
    .io_valid_29(InstBoard_io_valid_29),
    .io_valid_30(InstBoard_io_valid_30),
    .io_valid_31(InstBoard_io_valid_31),
    .io_RInstNo_1(InstBoard_io_RInstNo_1),
    .io_RInstNo_2(InstBoard_io_RInstNo_2),
    .io_RInstNo_3(InstBoard_io_RInstNo_3),
    .io_RInstNo_4(InstBoard_io_RInstNo_4),
    .io_RInstNo_5(InstBoard_io_RInstNo_5),
    .io_RInstNo_6(InstBoard_io_RInstNo_6),
    .io_RInstNo_7(InstBoard_io_RInstNo_7),
    .io_RInstNo_8(InstBoard_io_RInstNo_8),
    .io_RInstNo_9(InstBoard_io_RInstNo_9),
    .io_RInstNo_10(InstBoard_io_RInstNo_10),
    .io_RInstNo_11(InstBoard_io_RInstNo_11),
    .io_RInstNo_12(InstBoard_io_RInstNo_12),
    .io_RInstNo_13(InstBoard_io_RInstNo_13),
    .io_RInstNo_14(InstBoard_io_RInstNo_14),
    .io_RInstNo_15(InstBoard_io_RInstNo_15),
    .io_RInstNo_16(InstBoard_io_RInstNo_16),
    .io_RInstNo_17(InstBoard_io_RInstNo_17),
    .io_RInstNo_18(InstBoard_io_RInstNo_18),
    .io_RInstNo_19(InstBoard_io_RInstNo_19),
    .io_RInstNo_20(InstBoard_io_RInstNo_20),
    .io_RInstNo_21(InstBoard_io_RInstNo_21),
    .io_RInstNo_22(InstBoard_io_RInstNo_22),
    .io_RInstNo_23(InstBoard_io_RInstNo_23),
    .io_RInstNo_24(InstBoard_io_RInstNo_24),
    .io_RInstNo_25(InstBoard_io_RInstNo_25),
    .io_RInstNo_26(InstBoard_io_RInstNo_26),
    .io_RInstNo_27(InstBoard_io_RInstNo_27),
    .io_RInstNo_28(InstBoard_io_RInstNo_28),
    .io_RInstNo_29(InstBoard_io_RInstNo_29),
    .io_RInstNo_30(InstBoard_io_RInstNo_30),
    .io_RInstNo_31(InstBoard_io_RInstNo_31),
    .io_flush(InstBoard_io_flush)
  );
  InstQueue q ( // @[SIMD_ISU.scala 164:19]
    .clock(q_clock),
    .reset(q_reset),
    .io_setnum(q_io_setnum),
    .io_clearnum(q_io_clearnum),
    .io_HeadPtr(q_io_HeadPtr),
    .io_TailPtr(q_io_TailPtr),
    .io_Flag(q_io_Flag),
    .io_flush(q_io_flush)
  );
  assign io_in_0_ready = FrontisClear_1 | _T_521; // @[SIMD_ISU.scala 222:38]
  assign io_in_1_ready = ~io_in_1_valid | _T_524; // @[SIMD_ISU.scala 226:42]
  assign io_out_0_valid = io_in_0_valid & src1Ready_0 & src2Ready_0 & src3Ready_0 & ~(_T_480 & q_io_TailPtr !=
    q_io_HeadPtr); // @[SIMD_ISU.scala 215:141]
  assign io_out_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_runahead_checkpoint_id = io_in_0_bits_cf_runahead_checkpoint_id; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_cf_instrType = io_in_0_bits_cf_instrType; // @[SIMD_ISU.scala 247:27]
  assign io_out_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_funct3 = io_in_0_bits_ctrl_funct3; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_func24 = io_in_0_bits_ctrl_func24; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_func23 = io_in_0_bits_ctrl_func23; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_ctrl_isBru = io_in_0_bits_ctrl_fuOpType[4]; // @[ALU.scala 69:31]
  assign io_out_0_bits_ctrl_isMou = io_in_0_bits_ctrl_isMou; // @[SIMD_ISU.scala 248:29]
  assign io_out_0_bits_data_src1 = _T_592 | _T_590; // @[Mux.scala 27:72]
  assign io_out_0_bits_data_src2 = _T_724 | _T_722; // @[Mux.scala 27:72]
  assign io_out_0_bits_data_src3 = _T_1103 | _T_1102; // @[Mux.scala 27:72]
  assign io_out_0_bits_data_imm = io_in_0_bits_data_imm; // @[SIMD_ISU.scala 246:34]
  assign io_out_0_bits_InstNo = _T_1171[4:0]; // @[SIMD_ISU.scala 278:31]
  assign io_out_0_bits_InstFlag = _T_1168 ? ~q_io_Flag : q_io_Flag; // @[SIMD_ISU.scala 279:38]
  assign io_out_1_valid = io_in_1_valid & src1Ready_1 & src2Ready_1 & src3Ready_1 & ~RAWinIssue_1 & ~FrontHasCsrMouOp_1
     & ~(_T_505 & ~FrontisClear_1); // @[SIMD_ISU.scala 217:183]
  assign io_out_1_bits_cf_instr = io_in_1_bits_cf_instr; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_pc = io_in_1_bits_cf_pc; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_pnpc = io_in_1_bits_cf_pnpc; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_exceptionVec_1 = io_in_1_bits_cf_exceptionVec_1; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_exceptionVec_2 = io_in_1_bits_cf_exceptionVec_2; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_exceptionVec_12 = io_in_1_bits_cf_exceptionVec_12; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_0 = io_in_1_bits_cf_intrVec_0; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_1 = io_in_1_bits_cf_intrVec_1; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_2 = io_in_1_bits_cf_intrVec_2; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_3 = io_in_1_bits_cf_intrVec_3; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_4 = io_in_1_bits_cf_intrVec_4; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_5 = io_in_1_bits_cf_intrVec_5; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_6 = io_in_1_bits_cf_intrVec_6; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_7 = io_in_1_bits_cf_intrVec_7; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_8 = io_in_1_bits_cf_intrVec_8; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_9 = io_in_1_bits_cf_intrVec_9; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_10 = io_in_1_bits_cf_intrVec_10; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_intrVec_11 = io_in_1_bits_cf_intrVec_11; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_brIdx = io_in_1_bits_cf_brIdx; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_crossPageIPFFix = io_in_1_bits_cf_crossPageIPFFix; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_runahead_checkpoint_id = io_in_1_bits_cf_runahead_checkpoint_id; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_cf_instrType = io_in_1_bits_cf_instrType; // @[SIMD_ISU.scala 247:27]
  assign io_out_1_bits_ctrl_fuType = io_in_1_bits_ctrl_fuType; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_fuOpType = io_in_1_bits_ctrl_fuOpType; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_funct3 = io_in_1_bits_ctrl_funct3; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_func24 = io_in_1_bits_ctrl_func24; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_func23 = io_in_1_bits_ctrl_func23; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_rfWen = io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_rfDest = io_in_1_bits_ctrl_rfDest; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_ctrl_isBru = io_in_1_bits_ctrl_fuOpType[4]; // @[ALU.scala 69:31]
  assign io_out_1_bits_ctrl_isMou = io_in_1_bits_ctrl_isMou; // @[SIMD_ISU.scala 248:29]
  assign io_out_1_bits_data_src1 = _T_660 | _T_658; // @[Mux.scala 27:72]
  assign io_out_1_bits_data_src2 = _T_788 | _T_786; // @[Mux.scala 27:72]
  assign io_out_1_bits_data_src3 = _T_1162 | _T_1161; // @[Mux.scala 27:72]
  assign io_out_1_bits_data_imm = io_in_1_bits_data_imm; // @[SIMD_ISU.scala 246:34]
  assign io_out_1_bits_InstNo = _T_1178[4:0]; // @[SIMD_ISU.scala 278:31]
  assign io_out_1_bits_InstFlag = _T_1175 ? ~q_io_Flag : q_io_Flag; // @[SIMD_ISU.scala 279:38]
  assign io_wb_rfSrc1_0 = io_in_0_bits_ctrl_rfSrc1; // @[SIMD_ISU.scala 171:{25,25}]
  assign io_wb_rfSrc1_1 = io_in_1_bits_ctrl_rfSrc1; // @[SIMD_ISU.scala 171:{25,25}]
  assign io_wb_rfSrc2_0 = io_in_0_bits_ctrl_rfSrc2; // @[SIMD_ISU.scala 172:{25,25}]
  assign io_wb_rfSrc2_1 = io_in_1_bits_ctrl_rfSrc2; // @[SIMD_ISU.scala 172:{25,25}]
  assign io_wb_rfSrc3_0 = io_in_0_bits_ctrl_rfSrc3; // @[SIMD_ISU.scala 173:25 258:43]
  assign io_wb_rfSrc3_1 = io_in_1_bits_ctrl_rfSrc3; // @[SIMD_ISU.scala 173:25 258:43]
  assign io_TailPtr = q_io_TailPtr; // @[SIMD_ISU.scala 281:16]
  assign InstBoard_clock = clock;
  assign InstBoard_reset = reset;
  assign InstBoard_io_Wen_1 = 5'h1 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_2 = 5'h2 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h2 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_3 = 5'h3 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h3 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_4 = 5'h4 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h4 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_5 = 5'h5 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h5 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_6 = 5'h6 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h6 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_7 = 5'h7 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h7 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_8 = 5'h8 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h8 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_9 = 5'h9 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h9 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_10 = 5'ha == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'ha ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_11 = 5'hb == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'hb ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_12 = 5'hc == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'hc ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_13 = 5'hd == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'hd ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_14 = 5'he == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'he ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_15 = 5'hf == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'hf ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_16 = 5'h10 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h10 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_17 = 5'h11 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h11 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_18 = 5'h12 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h12 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_19 = 5'h13 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h13 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_20 = 5'h14 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h14 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_21 = 5'h15 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h15 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_22 = 5'h16 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h16 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_23 = 5'h17 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h17 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_24 = 5'h18 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h18 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_25 = 5'h19 == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h19 ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_26 = 5'h1a == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1a ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_27 = 5'h1b == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1b ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_28 = 5'h1c == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1c ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_29 = 5'h1d == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1d ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_30 = 5'h1e == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1e ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_Wen_31 = 5'h1f == io_in_0_bits_ctrl_rfDest & _T_521 & io_in_0_bits_ctrl_rfWen | 5'h1f ==
    io_in_1_bits_ctrl_rfDest & _T_524 & io_in_1_bits_ctrl_rfWen; // @[SIMD_ISU.scala 283:153]
  assign InstBoard_io_clear_1 = _T_1801 | io_wb_rfWen_7 & 5'h1 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_1; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_2 = _T_1840 | io_wb_rfWen_7 & 5'h2 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_2; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_3 = _T_1879 | io_wb_rfWen_7 & 5'h3 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_3; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_4 = _T_1918 | io_wb_rfWen_7 & 5'h4 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_4; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_5 = _T_1957 | io_wb_rfWen_7 & 5'h5 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_5; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_6 = _T_1996 | io_wb_rfWen_7 & 5'h6 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_6; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_7 = _T_2035 | io_wb_rfWen_7 & 5'h7 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_7; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_8 = _T_2074 | io_wb_rfWen_7 & 5'h8 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_8; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_9 = _T_2113 | io_wb_rfWen_7 & 5'h9 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_9; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_10 = _T_2152 | io_wb_rfWen_7 & 5'ha == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_10; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_11 = _T_2191 | io_wb_rfWen_7 & 5'hb == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_11; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_12 = _T_2230 | io_wb_rfWen_7 & 5'hc == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_12; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_13 = _T_2269 | io_wb_rfWen_7 & 5'hd == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_13; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_14 = _T_2308 | io_wb_rfWen_7 & 5'he == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_14; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_15 = _T_2347 | io_wb_rfWen_7 & 5'hf == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_15; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_16 = _T_2386 | io_wb_rfWen_7 & 5'h10 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_16; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_17 = _T_2425 | io_wb_rfWen_7 & 5'h11 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_17; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_18 = _T_2464 | io_wb_rfWen_7 & 5'h12 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_18; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_19 = _T_2503 | io_wb_rfWen_7 & 5'h13 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_19; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_20 = _T_2542 | io_wb_rfWen_7 & 5'h14 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_20; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_21 = _T_2581 | io_wb_rfWen_7 & 5'h15 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_21; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_22 = _T_2620 | io_wb_rfWen_7 & 5'h16 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_22; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_23 = _T_2659 | io_wb_rfWen_7 & 5'h17 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_23; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_24 = _T_2698 | io_wb_rfWen_7 & 5'h18 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_24; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_25 = _T_2737 | io_wb_rfWen_7 & 5'h19 == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_25; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_26 = _T_2776 | io_wb_rfWen_7 & 5'h1a == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_26; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_27 = _T_2815 | io_wb_rfWen_7 & 5'h1b == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_27; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_28 = _T_2854 | io_wb_rfWen_7 & 5'h1c == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_28; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_29 = _T_2893 | io_wb_rfWen_7 & 5'h1d == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_29; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_30 = _T_2932 | io_wb_rfWen_7 & 5'h1e == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_30; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_clear_31 = _T_2971 | io_wb_rfWen_7 & 5'h1f == io_wb_rfDest_7 & io_wb_InstNo_7 ==
    InstBoard_io_RInstNo_31; // @[SIMD_ISU.scala 291:197]
  assign InstBoard_io_WInstNo_1 = _T_1197 ? io_out_1_bits_InstNo : _GEN_482; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_2 = _T_1206 ? io_out_1_bits_InstNo : _GEN_484; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_3 = _T_1215 ? io_out_1_bits_InstNo : _GEN_486; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_4 = _T_1224 ? io_out_1_bits_InstNo : _GEN_488; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_5 = _T_1233 ? io_out_1_bits_InstNo : _GEN_490; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_6 = _T_1242 ? io_out_1_bits_InstNo : _GEN_492; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_7 = _T_1251 ? io_out_1_bits_InstNo : _GEN_494; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_8 = _T_1260 ? io_out_1_bits_InstNo : _GEN_496; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_9 = _T_1269 ? io_out_1_bits_InstNo : _GEN_498; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_10 = _T_1278 ? io_out_1_bits_InstNo : _GEN_500; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_11 = _T_1287 ? io_out_1_bits_InstNo : _GEN_502; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_12 = _T_1296 ? io_out_1_bits_InstNo : _GEN_504; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_13 = _T_1305 ? io_out_1_bits_InstNo : _GEN_506; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_14 = _T_1314 ? io_out_1_bits_InstNo : _GEN_508; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_15 = _T_1323 ? io_out_1_bits_InstNo : _GEN_510; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_16 = _T_1332 ? io_out_1_bits_InstNo : _GEN_512; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_17 = _T_1341 ? io_out_1_bits_InstNo : _GEN_514; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_18 = _T_1350 ? io_out_1_bits_InstNo : _GEN_516; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_19 = _T_1359 ? io_out_1_bits_InstNo : _GEN_518; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_20 = _T_1368 ? io_out_1_bits_InstNo : _GEN_520; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_21 = _T_1377 ? io_out_1_bits_InstNo : _GEN_522; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_22 = _T_1386 ? io_out_1_bits_InstNo : _GEN_524; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_23 = _T_1395 ? io_out_1_bits_InstNo : _GEN_526; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_24 = _T_1404 ? io_out_1_bits_InstNo : _GEN_528; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_25 = _T_1413 ? io_out_1_bits_InstNo : _GEN_530; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_26 = _T_1422 ? io_out_1_bits_InstNo : _GEN_532; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_27 = _T_1431 ? io_out_1_bits_InstNo : _GEN_534; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_28 = _T_1440 ? io_out_1_bits_InstNo : _GEN_536; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_29 = _T_1449 ? io_out_1_bits_InstNo : _GEN_538; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_30 = _T_1458 ? io_out_1_bits_InstNo : _GEN_540; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_WInstNo_31 = _T_1467 ? io_out_1_bits_InstNo : _GEN_542; // @[SIMD_ISU.scala 287:116 288:73]
  assign InstBoard_io_flush = io_flush; // @[SIMD_ISU.scala 292:26]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_setnum = {{3'd0}, _T_1166}; // @[SIMD_ISU.scala 272:17]
  assign q_io_clearnum = io_num_enterwbu; // @[SIMD_ISU.scala 274:18]
  assign q_io_flush = io_flush; // @[SIMD_ISU.scala 273:17]
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input  [38:0] io_cfIn_pnpc,
  input  [3:0]  io_cfIn_brIdx,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input  [63:0] io_offset
);
  wire  isAdderSub = ~io_in_bits_func[6]; // @[ALU.scala 94:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_in_bits_src2 ^ _T_2; // @[ALU.scala 95:33]
  wire [64:0] _T_4 = io_in_bits_src1 + _T_3; // @[ALU.scala 95:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 95:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 95:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[ALU.scala 96:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 97:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 98:28]
  wire [63:0] _T_10 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_14 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {_T_14,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_17 = 7'h25 == io_in_bits_func ? _T_10 : io_in_bits_src1; // @[Mux.scala 80:57]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[Mux.scala 80:57]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[ALU.scala 104:18]
  wire [126:0] _GEN_4 = {{63'd0}, shsrc1}; // @[ALU.scala 106:33]
  wire [126:0] _T_23 = _GEN_4 << shamt; // @[ALU.scala 106:33]
  wire [63:0] _T_25 = {63'h0,slt}; // @[Cat.scala 30:58]
  wire [63:0] _T_26 = {63'h0,sltu}; // @[Cat.scala 30:58]
  wire [63:0] _T_27 = shsrc1 >> shamt; // @[ALU.scala 110:32]
  wire [63:0] _T_28 = io_in_bits_src1 | io_in_bits_src2; // @[ALU.scala 111:30]
  wire [63:0] _T_29 = io_in_bits_src1 & io_in_bits_src2; // @[ALU.scala 112:30]
  wire [63:0] _T_30 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[ALU.scala 113:32]
  wire [63:0] _T_32 = $signed(_T_30) >>> shamt; // @[ALU.scala 113:49]
  wire [64:0] _T_34 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _T_23[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_36 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _T_25} : _T_34; // @[Mux.scala 80:57]
  wire [64:0] _T_38 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _T_26} : _T_36; // @[Mux.scala 80:57]
  wire [64:0] _T_40 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _T_38; // @[Mux.scala 80:57]
  wire [64:0] _T_42 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _T_27} : _T_40; // @[Mux.scala 80:57]
  wire [64:0] _T_44 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _T_28} : _T_42; // @[Mux.scala 80:57]
  wire [64:0] _T_46 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _T_29} : _T_44; // @[Mux.scala 80:57]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _T_32} : _T_46; // @[Mux.scala 80:57]
  wire [31:0] _T_52 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,res[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _T_53} : res; // @[ALU.scala 116:19]
  wire  _T_55 = ~(|xorRes); // @[ALU.scala 119:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[ALU.scala 70:30]
  wire  isBru = io_in_bits_func[4]; // @[ALU.scala 69:31]
  wire  _T_58 = 2'h0 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_59 = 2'h2 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = 2'h3 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_65 = _T_58 & _T_55 | _T_59 & slt | _T_60 & sltu; // @[Mux.scala 27:72]
  wire  taken = _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 126:72]
  wire [63:0] _GEN_1 = {{25'd0}, io_cfIn_pc}; // @[ALU.scala 127:41]
  wire [63:0] _T_68 = _GEN_1 + io_offset; // @[ALU.scala 127:41]
  wire [64:0] _T_69 = isBranch ? {{1'd0}, _T_68} : adderRes; // @[ALU.scala 127:19]
  wire [38:0] target = _T_69[38:0]; // @[ALU.scala 127:63]
  wire  _T_71 = ~taken & isBranch; // @[ALU.scala 128:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[ALU.scala 128:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 129:35]
  wire  _T_88 = ~isRVC; // @[ALU.scala 131:55]
  wire [38:0] _T_101 = io_cfIn_pc + 39'h2; // @[ALU.scala 132:71]
  wire [38:0] _T_103 = io_cfIn_pc + 39'h4; // @[ALU.scala 132:89]
  wire [38:0] _T_104 = isRVC ? _T_101 : _T_103; // @[ALU.scala 132:52]
  wire [24:0] _T_111 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_112 = {_T_111,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_114 = _T_112 + 64'h4; // @[ALU.scala 140:71]
  wire [63:0] _T_120 = _T_112 + 64'h2; // @[ALU.scala 140:108]
  wire [63:0] _T_121 = _T_88 ? _T_114 : _T_120; // @[ALU.scala 140:32]
  wire [64:0] _T_122 = isBru ? {{1'd0}, _T_121} : aluRes; // @[ALU.scala 140:21]
  assign io_out_bits = _T_122[63:0]; // @[ALU.scala 140:15]
  assign io_redirect_target = _T_71 ? _T_104 : target; // @[ALU.scala 132:28]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[ALU.scala 134:39]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:130 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 130:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fatal; // @[ALU.scala 130:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ALU_1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input  [38:0] io_cfIn_pnpc,
  input  [3:0]  io_cfIn_brIdx,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input  [63:0] io_offset
);
  wire  isAdderSub = ~io_in_bits_func[6]; // @[ALU.scala 94:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_in_bits_src2 ^ _T_2; // @[ALU.scala 95:33]
  wire [64:0] _T_4 = io_in_bits_src1 + _T_3; // @[ALU.scala 95:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 95:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 95:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[ALU.scala 96:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 97:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 98:28]
  wire [63:0] _T_10 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_14 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {_T_14,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_17 = 7'h25 == io_in_bits_func ? _T_10 : io_in_bits_src1; // @[Mux.scala 80:57]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[Mux.scala 80:57]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[ALU.scala 104:18]
  wire [126:0] _GEN_4 = {{63'd0}, shsrc1}; // @[ALU.scala 106:33]
  wire [126:0] _T_23 = _GEN_4 << shamt; // @[ALU.scala 106:33]
  wire [63:0] _T_25 = {63'h0,slt}; // @[Cat.scala 30:58]
  wire [63:0] _T_26 = {63'h0,sltu}; // @[Cat.scala 30:58]
  wire [63:0] _T_27 = shsrc1 >> shamt; // @[ALU.scala 110:32]
  wire [63:0] _T_28 = io_in_bits_src1 | io_in_bits_src2; // @[ALU.scala 111:30]
  wire [63:0] _T_29 = io_in_bits_src1 & io_in_bits_src2; // @[ALU.scala 112:30]
  wire [63:0] _T_30 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[ALU.scala 113:32]
  wire [63:0] _T_32 = $signed(_T_30) >>> shamt; // @[ALU.scala 113:49]
  wire [64:0] _T_34 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _T_23[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_36 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _T_25} : _T_34; // @[Mux.scala 80:57]
  wire [64:0] _T_38 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _T_26} : _T_36; // @[Mux.scala 80:57]
  wire [64:0] _T_40 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _T_38; // @[Mux.scala 80:57]
  wire [64:0] _T_42 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _T_27} : _T_40; // @[Mux.scala 80:57]
  wire [64:0] _T_44 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _T_28} : _T_42; // @[Mux.scala 80:57]
  wire [64:0] _T_46 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _T_29} : _T_44; // @[Mux.scala 80:57]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _T_32} : _T_46; // @[Mux.scala 80:57]
  wire [31:0] _T_52 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,res[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _T_53} : res; // @[ALU.scala 116:19]
  wire  _T_55 = ~(|xorRes); // @[ALU.scala 119:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[ALU.scala 70:30]
  wire  isBru = io_in_bits_func[4]; // @[ALU.scala 69:31]
  wire  _T_58 = 2'h0 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_59 = 2'h2 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = 2'h3 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_65 = _T_58 & _T_55 | _T_59 & slt | _T_60 & sltu; // @[Mux.scala 27:72]
  wire  taken = _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 126:72]
  wire [63:0] _GEN_1 = {{25'd0}, io_cfIn_pc}; // @[ALU.scala 127:41]
  wire [63:0] _T_68 = _GEN_1 + io_offset; // @[ALU.scala 127:41]
  wire [64:0] _T_69 = isBranch ? {{1'd0}, _T_68} : adderRes; // @[ALU.scala 127:19]
  wire [38:0] target = _T_69[38:0]; // @[ALU.scala 127:63]
  wire  _T_71 = ~taken & isBranch; // @[ALU.scala 128:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[ALU.scala 128:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 129:35]
  wire  _T_88 = ~isRVC; // @[ALU.scala 131:55]
  wire [38:0] _T_101 = io_cfIn_pc + 39'h2; // @[ALU.scala 132:71]
  wire [38:0] _T_103 = io_cfIn_pc + 39'h4; // @[ALU.scala 132:89]
  wire [38:0] _T_104 = isRVC ? _T_101 : _T_103; // @[ALU.scala 132:52]
  wire [24:0] _T_111 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_112 = {_T_111,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_114 = _T_112 + 64'h4; // @[ALU.scala 140:71]
  wire [63:0] _T_120 = _T_112 + 64'h2; // @[ALU.scala 140:108]
  wire [63:0] _T_121 = _T_88 ? _T_114 : _T_120; // @[ALU.scala 140:32]
  wire [64:0] _T_122 = isBru ? {{1'd0}, _T_121} : aluRes; // @[ALU.scala 140:21]
  assign io_out_bits = _T_122[63:0]; // @[ALU.scala 140:15]
  assign io_redirect_target = _T_71 ? _T_104 : target; // @[ALU.scala 132:28]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[ALU.scala 134:39]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:130 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 130:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fatal; // @[ALU.scala 130:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PALU(
  output        io_in_ready,
  input         io_in_valid,
  input  [38:0] io_in_bits_DecodeIn_cf_pc,
  input  [63:0] io_in_bits_DecodeIn_cf_runahead_checkpoint_id,
  input  [6:0]  io_in_bits_DecodeIn_ctrl_fuOpType,
  input  [2:0]  io_in_bits_DecodeIn_ctrl_funct3,
  input         io_in_bits_DecodeIn_ctrl_func24,
  input         io_in_bits_DecodeIn_ctrl_rfWen,
  input  [4:0]  io_in_bits_DecodeIn_ctrl_rfDest,
  input  [63:0] io_in_bits_DecodeIn_data_src1,
  input  [63:0] io_in_bits_DecodeIn_data_src2,
  input  [63:0] io_in_bits_DecodeIn_data_src3,
  input  [4:0]  io_in_bits_DecodeIn_InstNo,
  input         io_in_bits_DecodeIn_InstFlag,
  input         io_in_bits_Pctrl_isAdd_64,
  input         io_in_bits_Pctrl_isAdd_32,
  input         io_in_bits_Pctrl_isAdd_16,
  input         io_in_bits_Pctrl_isAdd_8,
  input         io_in_bits_Pctrl_isAdd_Q15,
  input         io_in_bits_Pctrl_isAdd_Q31,
  input         io_in_bits_Pctrl_isAdd_C31,
  input         io_in_bits_Pctrl_isAve,
  input         io_in_bits_Pctrl_isSub_64,
  input         io_in_bits_Pctrl_isSub_32,
  input         io_in_bits_Pctrl_isSub_16,
  input         io_in_bits_Pctrl_isSub_8,
  input         io_in_bits_Pctrl_isSub_Q15,
  input         io_in_bits_Pctrl_isSub_Q31,
  input         io_in_bits_Pctrl_isSub_C31,
  input         io_in_bits_Pctrl_isCras_16,
  input         io_in_bits_Pctrl_isCrsa_16,
  input         io_in_bits_Pctrl_isCras_32,
  input         io_in_bits_Pctrl_isCrsa_32,
  input         io_in_bits_Pctrl_isStas_16,
  input         io_in_bits_Pctrl_isStsa_16,
  input         io_in_bits_Pctrl_isStas_32,
  input         io_in_bits_Pctrl_isStsa_32,
  input         io_in_bits_Pctrl_isComp_16,
  input         io_in_bits_Pctrl_isComp_8,
  input         io_in_bits_Pctrl_isCompare,
  input         io_in_bits_Pctrl_isMaxMin_16,
  input         io_in_bits_Pctrl_isMaxMin_8,
  input         io_in_bits_Pctrl_isMaxMin_XLEN,
  input         io_in_bits_Pctrl_isMaxMin_32,
  input         io_in_bits_Pctrl_isMaxMin,
  input         io_in_bits_Pctrl_isPbs,
  input         io_in_bits_Pctrl_isRs_16,
  input         io_in_bits_Pctrl_isLs_16,
  input         io_in_bits_Pctrl_isLR_16,
  input         io_in_bits_Pctrl_isRs_8,
  input         io_in_bits_Pctrl_isLs_8,
  input         io_in_bits_Pctrl_isLR_8,
  input         io_in_bits_Pctrl_isRs_32,
  input         io_in_bits_Pctrl_isLs_32,
  input         io_in_bits_Pctrl_isLR_32,
  input         io_in_bits_Pctrl_isLR_Q31,
  input         io_in_bits_Pctrl_isLs_Q31,
  input         io_in_bits_Pctrl_isRs_XLEN,
  input         io_in_bits_Pctrl_isSRAIWU,
  input         io_in_bits_Pctrl_isFSRW,
  input         io_in_bits_Pctrl_isWext,
  input         io_in_bits_Pctrl_isShifter,
  input         io_in_bits_Pctrl_isClip_16,
  input         io_in_bits_Pctrl_isClip_8,
  input         io_in_bits_Pctrl_isclip_32,
  input         io_in_bits_Pctrl_isClip,
  input         io_in_bits_Pctrl_isSat_16,
  input         io_in_bits_Pctrl_isSat_8,
  input         io_in_bits_Pctrl_isSat_32,
  input         io_in_bits_Pctrl_isSat_W,
  input         io_in_bits_Pctrl_isSat,
  input         io_in_bits_Pctrl_isCnt_16,
  input         io_in_bits_Pctrl_isCnt_8,
  input         io_in_bits_Pctrl_isCnt_32,
  input         io_in_bits_Pctrl_isCnt,
  input         io_in_bits_Pctrl_isSwap_16,
  input         io_in_bits_Pctrl_isSwap_8,
  input         io_in_bits_Pctrl_isSwap,
  input         io_in_bits_Pctrl_isUnpack,
  input         io_in_bits_Pctrl_isBitrev,
  input         io_in_bits_Pctrl_isCmix,
  input         io_in_bits_Pctrl_isInsertb,
  input         io_in_bits_Pctrl_isPackbb,
  input         io_in_bits_Pctrl_isPackbt,
  input         io_in_bits_Pctrl_isPacktb,
  input         io_in_bits_Pctrl_isPacktt,
  input         io_in_bits_Pctrl_isPack,
  input  [7:0]  io_in_bits_Pctrl_isSub,
  input         io_in_bits_Pctrl_isAdder,
  input         io_in_bits_Pctrl_SrcSigned,
  input         io_in_bits_Pctrl_Saturating,
  input         io_in_bits_Pctrl_Translation,
  input         io_in_bits_Pctrl_LessEqual,
  input         io_in_bits_Pctrl_LessThan,
  input  [79:0] io_in_bits_Pctrl_adderRes_ori,
  input  [63:0] io_in_bits_Pctrl_adderRes,
  input  [79:0] io_in_bits_Pctrl_adderRes_ori_drophighestbit,
  input         io_in_bits_Pctrl_Round,
  input         io_in_bits_Pctrl_ShiftSigned,
  input         io_in_bits_Pctrl_Arithmetic,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_result,
  output [38:0] io_out_bits_DecodeOut_cf_pc,
  output [63:0] io_out_bits_DecodeOut_cf_runahead_checkpoint_id,
  output        io_out_bits_DecodeOut_ctrl_rfWen,
  output [4:0]  io_out_bits_DecodeOut_ctrl_rfDest,
  output        io_out_bits_DecodeOut_pext_OV,
  output [4:0]  io_out_bits_DecodeOut_InstNo,
  output        io_out_bits_DecodeOut_InstFlag
);
  wire  _T_1 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15; // @[PALU.scala 186:43]
  wire  _T_15 = ~io_in_bits_DecodeIn_ctrl_fuOpType[3]; // @[PALU.scala 186:55]
  wire  _T_16 = io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15 ? ~io_in_bits_DecodeIn_ctrl_fuOpType[3] :
    io_in_bits_Pctrl_SrcSigned; // @[PALU.scala 186:33]
  wire  _GEN_7 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[17] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[15] :
    io_in_bits_Pctrl_adderRes_ori[16]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_0 = io_in_bits_Pctrl_adderRes_ori[17] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_1 = _GEN_7 ? _GEN_0 : io_in_bits_Pctrl_adderRes_ori[15:0]; // @[PALU.scala 123:21 126:33]
  wire [15:0] _GEN_3 = io_in_bits_Pctrl_isSub[0] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_5 = _GEN_7 ? _GEN_3 : io_in_bits_Pctrl_adderRes_ori[15:0]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_8 = _T_16 ? _GEN_1 : _GEN_5; // @[PALU.scala 124:28]
  wire  _GEN_17 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[35] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[33] :
    io_in_bits_Pctrl_adderRes_ori[34]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_10 = io_in_bits_Pctrl_adderRes_ori[35] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_11 = _GEN_17 ? _GEN_10 : io_in_bits_Pctrl_adderRes_ori[33:18]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_12 = _GEN_17 | _GEN_7; // @[PALU.scala 126:33 132:24]
  wire [15:0] _GEN_13 = io_in_bits_Pctrl_isSub[1] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_15 = _GEN_17 ? _GEN_13 : io_in_bits_Pctrl_adderRes_ori[33:18]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_18 = _T_16 ? _GEN_11 : _GEN_15; // @[PALU.scala 124:28]
  wire  _GEN_19 = _T_16 ? _GEN_12 : _GEN_12; // @[PALU.scala 124:28]
  wire  _GEN_27 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[53] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[51] :
    io_in_bits_Pctrl_adderRes_ori[52]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_20 = io_in_bits_Pctrl_adderRes_ori[53] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_21 = _GEN_27 ? _GEN_20 : io_in_bits_Pctrl_adderRes_ori[51:36]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_22 = _GEN_27 | _GEN_19; // @[PALU.scala 126:33 132:24]
  wire [15:0] _GEN_23 = io_in_bits_Pctrl_isSub[2] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_25 = _GEN_27 ? _GEN_23 : io_in_bits_Pctrl_adderRes_ori[51:36]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_28 = _T_16 ? _GEN_21 : _GEN_25; // @[PALU.scala 124:28]
  wire  _GEN_29 = _T_16 ? _GEN_22 : _GEN_22; // @[PALU.scala 124:28]
  wire  _GEN_37 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[71] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[69] :
    io_in_bits_Pctrl_adderRes_ori[70]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_30 = io_in_bits_Pctrl_adderRes_ori[71] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_31 = _GEN_37 ? _GEN_30 : io_in_bits_Pctrl_adderRes_ori[69:54]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_32 = _GEN_37 | _GEN_29; // @[PALU.scala 126:33 132:24]
  wire [15:0] _GEN_33 = io_in_bits_Pctrl_isSub[3] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_35 = _GEN_37 ? _GEN_33 : io_in_bits_Pctrl_adderRes_ori[69:54]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_38 = _T_16 ? _GEN_31 : _GEN_35; // @[PALU.scala 124:28]
  wire  _GEN_39 = _T_16 ? _GEN_32 : _GEN_32; // @[PALU.scala 124:28]
  wire [64:0] _T_80 = {_GEN_39,_GEN_38,_GEN_28,_GEN_18,_GEN_8}; // @[Cat.scala 30:58]
  wire [47:0] _T_85 = _T_80[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_86 = {_T_85,_T_80[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_88 = _T_12 ? _T_86 : _T_80[63:0]; // @[PALU.scala 188:34]
  wire [63:0] _T_101 = {io_in_bits_Pctrl_adderRes_ori[70:55],io_in_bits_Pctrl_adderRes_ori[52:37],
    io_in_bits_Pctrl_adderRes_ori[34:19],io_in_bits_Pctrl_adderRes_ori[16:1]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_40 = io_in_bits_Pctrl_Translation ? _T_101 : io_in_bits_Pctrl_adderRes; // @[PALU.scala 190:32 191:28]
  wire [63:0] _GEN_41 = io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15 ? _T_88 :
    _GEN_40; // @[PALU.scala 185:49 188:28]
  wire  _GEN_42 = (io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15) & _T_80[64]; // @[PALU.scala 185:49 189:21]
  wire  _GEN_50 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[9] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[7] : io_in_bits_Pctrl_adderRes_ori[8]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_43 = io_in_bits_Pctrl_adderRes_ori[9] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_44 = _GEN_50 ? _GEN_43 : io_in_bits_Pctrl_adderRes_ori[7:0]; // @[PALU.scala 123:21 126:33]
  wire [7:0] _GEN_46 = io_in_bits_Pctrl_isSub[0] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_48 = _GEN_50 ? _GEN_46 : io_in_bits_Pctrl_adderRes_ori[7:0]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_51 = io_in_bits_Pctrl_SrcSigned ? _GEN_44 : _GEN_48; // @[PALU.scala 124:28]
  wire  _GEN_60 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[19] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[17] : io_in_bits_Pctrl_adderRes_ori[18]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_53 = io_in_bits_Pctrl_adderRes_ori[19] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_54 = _GEN_60 ? _GEN_53 : io_in_bits_Pctrl_adderRes_ori[17:10]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_55 = _GEN_60 | _GEN_50; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_56 = io_in_bits_Pctrl_isSub[1] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_58 = _GEN_60 ? _GEN_56 : io_in_bits_Pctrl_adderRes_ori[17:10]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_61 = io_in_bits_Pctrl_SrcSigned ? _GEN_54 : _GEN_58; // @[PALU.scala 124:28]
  wire  _GEN_62 = io_in_bits_Pctrl_SrcSigned ? _GEN_55 : _GEN_55; // @[PALU.scala 124:28]
  wire  _GEN_70 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[29] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[27] : io_in_bits_Pctrl_adderRes_ori[28]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_63 = io_in_bits_Pctrl_adderRes_ori[29] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_64 = _GEN_70 ? _GEN_63 : io_in_bits_Pctrl_adderRes_ori[27:20]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_65 = _GEN_70 | _GEN_62; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_66 = io_in_bits_Pctrl_isSub[2] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_68 = _GEN_70 ? _GEN_66 : io_in_bits_Pctrl_adderRes_ori[27:20]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_71 = io_in_bits_Pctrl_SrcSigned ? _GEN_64 : _GEN_68; // @[PALU.scala 124:28]
  wire  _GEN_72 = io_in_bits_Pctrl_SrcSigned ? _GEN_65 : _GEN_65; // @[PALU.scala 124:28]
  wire  _GEN_80 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[39] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[37] : io_in_bits_Pctrl_adderRes_ori[38]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_73 = io_in_bits_Pctrl_adderRes_ori[39] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_74 = _GEN_80 ? _GEN_73 : io_in_bits_Pctrl_adderRes_ori[37:30]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_75 = _GEN_80 | _GEN_72; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_76 = io_in_bits_Pctrl_isSub[3] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_78 = _GEN_80 ? _GEN_76 : io_in_bits_Pctrl_adderRes_ori[37:30]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_81 = io_in_bits_Pctrl_SrcSigned ? _GEN_74 : _GEN_78; // @[PALU.scala 124:28]
  wire  _GEN_82 = io_in_bits_Pctrl_SrcSigned ? _GEN_75 : _GEN_75; // @[PALU.scala 124:28]
  wire  _GEN_90 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[49] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[47] : io_in_bits_Pctrl_adderRes_ori[48]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_83 = io_in_bits_Pctrl_adderRes_ori[49] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_84 = _GEN_90 ? _GEN_83 : io_in_bits_Pctrl_adderRes_ori[47:40]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_85 = _GEN_90 | _GEN_82; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_86 = io_in_bits_Pctrl_isSub[4] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_88 = _GEN_90 ? _GEN_86 : io_in_bits_Pctrl_adderRes_ori[47:40]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_91 = io_in_bits_Pctrl_SrcSigned ? _GEN_84 : _GEN_88; // @[PALU.scala 124:28]
  wire  _GEN_92 = io_in_bits_Pctrl_SrcSigned ? _GEN_85 : _GEN_85; // @[PALU.scala 124:28]
  wire  _GEN_100 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[59] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[57] : io_in_bits_Pctrl_adderRes_ori[58]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_93 = io_in_bits_Pctrl_adderRes_ori[59] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_94 = _GEN_100 ? _GEN_93 : io_in_bits_Pctrl_adderRes_ori[57:50]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_95 = _GEN_100 | _GEN_92; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_96 = io_in_bits_Pctrl_isSub[5] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_98 = _GEN_100 ? _GEN_96 : io_in_bits_Pctrl_adderRes_ori[57:50]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_101 = io_in_bits_Pctrl_SrcSigned ? _GEN_94 : _GEN_98; // @[PALU.scala 124:28]
  wire  _GEN_102 = io_in_bits_Pctrl_SrcSigned ? _GEN_95 : _GEN_95; // @[PALU.scala 124:28]
  wire  _GEN_110 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[69] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[67] : io_in_bits_Pctrl_adderRes_ori[68]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_103 = io_in_bits_Pctrl_adderRes_ori[69] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_104 = _GEN_110 ? _GEN_103 : io_in_bits_Pctrl_adderRes_ori[67:60]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_105 = _GEN_110 | _GEN_102; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_106 = io_in_bits_Pctrl_isSub[6] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_108 = _GEN_110 ? _GEN_106 : io_in_bits_Pctrl_adderRes_ori[67:60]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_111 = io_in_bits_Pctrl_SrcSigned ? _GEN_104 : _GEN_108; // @[PALU.scala 124:28]
  wire  _GEN_112 = io_in_bits_Pctrl_SrcSigned ? _GEN_105 : _GEN_105; // @[PALU.scala 124:28]
  wire  _GEN_120 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[79] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[77] : io_in_bits_Pctrl_adderRes_ori[78]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_113 = io_in_bits_Pctrl_adderRes_ori[79] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_114 = _GEN_120 ? _GEN_113 : io_in_bits_Pctrl_adderRes_ori[77:70]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_115 = _GEN_120 | _GEN_112; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_116 = io_in_bits_Pctrl_isSub[7] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_118 = _GEN_120 ? _GEN_116 : io_in_bits_Pctrl_adderRes_ori[77:70]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_121 = io_in_bits_Pctrl_SrcSigned ? _GEN_114 : _GEN_118; // @[PALU.scala 124:28]
  wire  _GEN_122 = io_in_bits_Pctrl_SrcSigned ? _GEN_115 : _GEN_115; // @[PALU.scala 124:28]
  wire [64:0] _T_230 = {_GEN_122,_GEN_121,_GEN_111,_GEN_101,_GEN_91,_GEN_81,_GEN_71,_GEN_61,_GEN_51}; // @[Cat.scala 30:58]
  wire [63:0] _T_256 = {io_in_bits_Pctrl_adderRes_ori[78:71],io_in_bits_Pctrl_adderRes_ori[68:61],
    io_in_bits_Pctrl_adderRes_ori[58:51],io_in_bits_Pctrl_adderRes_ori[48:41],io_in_bits_Pctrl_adderRes_ori[38:31],
    io_in_bits_Pctrl_adderRes_ori[28:21],io_in_bits_Pctrl_adderRes_ori[18:11],io_in_bits_Pctrl_adderRes_ori[8:1]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_123 = io_in_bits_Pctrl_Translation ? _T_256 : io_in_bits_Pctrl_adderRes; // @[PALU.scala 198:32 199:28]
  wire [63:0] _GEN_124 = io_in_bits_Pctrl_Saturating ? _T_230[63:0] : _GEN_123; // @[PALU.scala 194:25 196:28]
  wire  _GEN_125 = io_in_bits_Pctrl_Saturating & _T_230[64]; // @[PALU.scala 194:25 197:21]
  wire  _T_266 = io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31; // @[PALU.scala 203:44]
  wire  _T_270 = io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31 ? _T_15 : io_in_bits_Pctrl_SrcSigned; // @[PALU.scala 203:33]
  wire  _GEN_133 = _T_270 ? io_in_bits_Pctrl_adderRes_ori[33] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[31] :
    io_in_bits_Pctrl_adderRes_ori[32]; // @[PALU.scala 124:28 125:21 135:21]
  wire [31:0] _GEN_126 = io_in_bits_Pctrl_adderRes_ori[33] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 127:66 128:33 130:33]
  wire [31:0] _GEN_127 = _GEN_133 ? _GEN_126 : io_in_bits_Pctrl_adderRes_ori[31:0]; // @[PALU.scala 123:21 126:33]
  wire [31:0] _GEN_129 = io_in_bits_Pctrl_isSub[0] ? 32'h0 : 32'hffffffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [31:0] _GEN_131 = _GEN_133 ? _GEN_129 : io_in_bits_Pctrl_adderRes_ori[31:0]; // @[PALU.scala 123:21 136:33]
  wire [31:0] _GEN_134 = _T_270 ? _GEN_127 : _GEN_131; // @[PALU.scala 124:28]
  wire  _GEN_143 = _T_270 ? io_in_bits_Pctrl_adderRes_ori[67] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[65] :
    io_in_bits_Pctrl_adderRes_ori[66]; // @[PALU.scala 124:28 125:21 135:21]
  wire [31:0] _GEN_136 = io_in_bits_Pctrl_adderRes_ori[67] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 127:66 128:33 130:33]
  wire [31:0] _GEN_137 = _GEN_143 ? _GEN_136 : io_in_bits_Pctrl_adderRes_ori[65:34]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_138 = _GEN_143 | _GEN_133; // @[PALU.scala 126:33 132:24]
  wire [31:0] _GEN_139 = io_in_bits_Pctrl_isSub[1] ? 32'h0 : 32'hffffffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [31:0] _GEN_141 = _GEN_143 ? _GEN_139 : io_in_bits_Pctrl_adderRes_ori[65:34]; // @[PALU.scala 123:21 136:33]
  wire [31:0] _GEN_144 = _T_270 ? _GEN_137 : _GEN_141; // @[PALU.scala 124:28]
  wire  _GEN_145 = _T_270 ? _GEN_138 : _GEN_138; // @[PALU.scala 124:28]
  wire [64:0] _T_302 = {_GEN_145,_GEN_144,_GEN_134}; // @[Cat.scala 30:58]
  wire [31:0] _T_307 = _T_302[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_308 = {_T_307,_T_302[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_310 = _T_266 ? _T_308 : _T_302[63:0]; // @[PALU.scala 205:34]
  wire [63:0] _T_317 = {io_in_bits_Pctrl_adderRes_ori[66:35],io_in_bits_Pctrl_adderRes_ori[32:1]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_146 = io_in_bits_Pctrl_Translation ? _T_317 : io_in_bits_Pctrl_adderRes; // @[PALU.scala 207:32 208:28]
  wire [63:0] _GEN_147 = io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31 ? _T_310
     : _GEN_146; // @[PALU.scala 202:49 205:28]
  wire  _GEN_148 = (io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31) & _T_302[64]; // @[PALU.scala 202:49 206:21]
  wire  _GEN_156 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[65] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[63] : io_in_bits_Pctrl_adderRes_ori[64]; // @[PALU.scala 124:28 125:21 135:21]
  wire [63:0] _GEN_149 = io_in_bits_Pctrl_adderRes_ori[65] ? 64'h8000000000000000 : 64'h7fffffffffffffff; // @[PALU.scala 127:66 128:33 130:33]
  wire [63:0] _GEN_150 = _GEN_156 ? _GEN_149 : io_in_bits_Pctrl_adderRes_ori[63:0]; // @[PALU.scala 123:21 126:33]
  wire [63:0] _GEN_152 = io_in_bits_Pctrl_isSub[0] ? 64'h0 : 64'hffffffffffffffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [63:0] _GEN_154 = _GEN_156 ? _GEN_152 : io_in_bits_Pctrl_adderRes_ori[63:0]; // @[PALU.scala 123:21 136:33]
  wire [63:0] _GEN_157 = io_in_bits_Pctrl_SrcSigned ? _GEN_150 : _GEN_154; // @[PALU.scala 124:28]
  wire [64:0] _T_334 = {_GEN_156,_GEN_157}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_159 = io_in_bits_Pctrl_Translation ? io_in_bits_Pctrl_adderRes_ori[64:1] : io_in_bits_Pctrl_adderRes; // @[PALU.scala 215:32 216:28]
  wire [63:0] _GEN_160 = io_in_bits_Pctrl_Saturating ? _T_334[63:0] : _GEN_159; // @[PALU.scala 211:25 213:28]
  wire  _GEN_161 = io_in_bits_Pctrl_Saturating & _T_334[64]; // @[PALU.scala 211:25 214:21]
  wire [31:0] _T_349 = _T_317[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_350 = {_T_349,_T_317[31:0]}; // @[Cat.scala 30:58]
  wire [80:0] _T_351 = io_in_bits_Pctrl_adderRes_ori + 80'h1; // @[PALU.scala 221:40]
  wire [63:0] _GEN_162 = io_in_bits_Pctrl_isAve ? _T_351[64:1] : io_in_bits_Pctrl_adderRes; // @[PALU.scala 220:22 221:24]
  wire [63:0] _GEN_163 = io_in_bits_Pctrl_isSub_C31 | io_in_bits_Pctrl_isAdd_C31 ? _T_350 : _GEN_162; // @[PALU.scala 218:37 219:24]
  wire [63:0] _GEN_164 = io_in_bits_Pctrl_isAdd_64 | io_in_bits_Pctrl_isSub_64 ? _GEN_160 : _GEN_163; // @[PALU.scala 210:36]
  wire  _GEN_165 = (io_in_bits_Pctrl_isAdd_64 | io_in_bits_Pctrl_isSub_64) & _GEN_161; // @[PALU.scala 210:36]
  wire [63:0] _GEN_166 = io_in_bits_Pctrl_isAdd_32 | io_in_bits_Pctrl_isSub_32 | io_in_bits_Pctrl_isCras_32 |
    io_in_bits_Pctrl_isCrsa_32 | io_in_bits_Pctrl_isStas_32 | io_in_bits_Pctrl_isStsa_32 | io_in_bits_Pctrl_isAdd_Q31 |
    io_in_bits_Pctrl_isSub_Q31 ? _GEN_147 : _GEN_164; // @[PALU.scala 201:108]
  wire  _GEN_167 = io_in_bits_Pctrl_isAdd_32 | io_in_bits_Pctrl_isSub_32 | io_in_bits_Pctrl_isCras_32 |
    io_in_bits_Pctrl_isCrsa_32 | io_in_bits_Pctrl_isStas_32 | io_in_bits_Pctrl_isStsa_32 | io_in_bits_Pctrl_isAdd_Q31 |
    io_in_bits_Pctrl_isSub_Q31 ? _GEN_148 : _GEN_165; // @[PALU.scala 201:108]
  wire [63:0] _GEN_168 = io_in_bits_Pctrl_isAdd_8 | io_in_bits_Pctrl_isSub_8 ? _GEN_124 : _GEN_166; // @[PALU.scala 193:34]
  wire  _GEN_169 = io_in_bits_Pctrl_isAdd_8 | io_in_bits_Pctrl_isSub_8 ? _GEN_125 : _GEN_167; // @[PALU.scala 193:34]
  wire [63:0] adderRes_final = io_in_bits_Pctrl_isAdd_16 | io_in_bits_Pctrl_isSub_16 | io_in_bits_Pctrl_isCras_16 |
    io_in_bits_Pctrl_isCrsa_16 | io_in_bits_Pctrl_isStas_16 | io_in_bits_Pctrl_isStsa_16 | io_in_bits_Pctrl_isAdd_Q15 |
    io_in_bits_Pctrl_isSub_Q15 ? _GEN_41 : _GEN_168; // @[PALU.scala 184:101]
  wire  adderOV = io_in_bits_Pctrl_isAdd_16 | io_in_bits_Pctrl_isSub_16 | io_in_bits_Pctrl_isCras_16 |
    io_in_bits_Pctrl_isCrsa_16 | io_in_bits_Pctrl_isStas_16 | io_in_bits_Pctrl_isStsa_16 | io_in_bits_Pctrl_isAdd_Q15 |
    io_in_bits_Pctrl_isSub_Q15 ? _GEN_42 : _GEN_169; // @[PALU.scala 184:101]
  wire  _T_356 = io_in_bits_Pctrl_adderRes_ori[15:0] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_358 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[16] | _T_356 : _T_356; // @[PALU.scala 164:55]
  wire  _T_359 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[16] : _T_358; // @[PALU.scala 164:31]
  wire [15:0] _T_361 = _T_359 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire  _T_365 = io_in_bits_Pctrl_adderRes_ori[33:18] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_367 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[34] | _T_365 : _T_365; // @[PALU.scala 164:55]
  wire  _T_368 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[34] : _T_367; // @[PALU.scala 164:31]
  wire [15:0] _T_370 = _T_368 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire  _T_374 = io_in_bits_Pctrl_adderRes_ori[51:36] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_376 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[52] | _T_374 : _T_374; // @[PALU.scala 164:55]
  wire  _T_377 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[52] : _T_376; // @[PALU.scala 164:31]
  wire [15:0] _T_379 = _T_377 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire  _T_383 = io_in_bits_Pctrl_adderRes_ori[69:54] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_385 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[70] | _T_383 : _T_383; // @[PALU.scala 164:55]
  wire  _T_386 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[70] : _T_385; // @[PALU.scala 164:31]
  wire [15:0] _T_388 = _T_386 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_391 = {_T_388,_T_379,_T_370,_T_361}; // @[Cat.scala 30:58]
  wire  _T_395 = io_in_bits_Pctrl_adderRes_ori[7:0] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_397 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[8] | _T_395 : _T_395; // @[PALU.scala 164:55]
  wire  _T_398 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[8] : _T_397; // @[PALU.scala 164:31]
  wire [7:0] _T_400 = _T_398 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_404 = io_in_bits_Pctrl_adderRes_ori[17:10] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_406 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[18] | _T_404 : _T_404; // @[PALU.scala 164:55]
  wire  _T_407 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[18] : _T_406; // @[PALU.scala 164:31]
  wire [7:0] _T_409 = _T_407 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_413 = io_in_bits_Pctrl_adderRes_ori[27:20] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_415 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[28] | _T_413 : _T_413; // @[PALU.scala 164:55]
  wire  _T_416 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[28] : _T_415; // @[PALU.scala 164:31]
  wire [7:0] _T_418 = _T_416 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_422 = io_in_bits_Pctrl_adderRes_ori[37:30] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_424 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[38] | _T_422 : _T_422; // @[PALU.scala 164:55]
  wire  _T_425 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[38] : _T_424; // @[PALU.scala 164:31]
  wire [7:0] _T_427 = _T_425 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_431 = io_in_bits_Pctrl_adderRes_ori[47:40] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_433 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[48] | _T_431 : _T_431; // @[PALU.scala 164:55]
  wire  _T_434 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[48] : _T_433; // @[PALU.scala 164:31]
  wire [7:0] _T_436 = _T_434 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_440 = io_in_bits_Pctrl_adderRes_ori[57:50] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_442 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[58] | _T_440 : _T_440; // @[PALU.scala 164:55]
  wire  _T_443 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[58] : _T_442; // @[PALU.scala 164:31]
  wire [7:0] _T_445 = _T_443 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_449 = io_in_bits_Pctrl_adderRes_ori[67:60] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_451 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[68] | _T_449 : _T_449; // @[PALU.scala 164:55]
  wire  _T_452 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[68] : _T_451; // @[PALU.scala 164:31]
  wire [7:0] _T_454 = _T_452 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_458 = io_in_bits_Pctrl_adderRes_ori[77:70] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_460 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[78] | _T_458 : _T_458; // @[PALU.scala 164:55]
  wire  _T_461 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[78] : _T_460; // @[PALU.scala 164:31]
  wire [7:0] _T_463 = _T_461 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_470 = {_T_463,_T_454,_T_445,_T_436,_T_427,_T_418,_T_409,_T_400}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_172 = io_in_bits_Pctrl_isComp_8 ? _T_470 : 64'h0; // @[PALU.scala 228:25 229:20]
  wire [63:0] compareRes = io_in_bits_Pctrl_isComp_16 ? _T_391 : _GEN_172; // @[PALU.scala 226:20 227:20]
  wire  _T_473 = ~io_in_bits_DecodeIn_ctrl_fuOpType[0]; // @[PALU.scala 235:55]
  wire [15:0] _T_480 = ~(io_in_bits_Pctrl_adderRes_ori[16] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[15:0] :
    io_in_bits_DecodeIn_data_src2[15:0]; // @[PALU.scala 175:30]
  wire [15:0] _T_498 = ~(io_in_bits_Pctrl_adderRes_ori[34] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[31:16] :
    io_in_bits_DecodeIn_data_src2[31:16]; // @[PALU.scala 175:30]
  wire [15:0] _T_516 = ~(io_in_bits_Pctrl_adderRes_ori[52] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[47:32] :
    io_in_bits_DecodeIn_data_src2[47:32]; // @[PALU.scala 175:30]
  wire [15:0] _T_534 = ~(io_in_bits_Pctrl_adderRes_ori[70] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[63:48] :
    io_in_bits_DecodeIn_data_src2[63:48]; // @[PALU.scala 175:30]
  wire [63:0] _T_548 = {_T_534,_T_516,_T_498,_T_480}; // @[Cat.scala 30:58]
  wire [7:0] _T_558 = ~(io_in_bits_Pctrl_adderRes_ori[8] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src2[7:0]; // @[PALU.scala 175:30]
  wire [7:0] _T_576 = ~(io_in_bits_Pctrl_adderRes_ori[18] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[15:8] :
    io_in_bits_DecodeIn_data_src2[15:8]; // @[PALU.scala 175:30]
  wire [7:0] _T_594 = ~(io_in_bits_Pctrl_adderRes_ori[28] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[23:16] :
    io_in_bits_DecodeIn_data_src2[23:16]; // @[PALU.scala 175:30]
  wire [7:0] _T_612 = ~(io_in_bits_Pctrl_adderRes_ori[38] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[31:24] :
    io_in_bits_DecodeIn_data_src2[31:24]; // @[PALU.scala 175:30]
  wire [7:0] _T_630 = ~(io_in_bits_Pctrl_adderRes_ori[48] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[39:32] :
    io_in_bits_DecodeIn_data_src2[39:32]; // @[PALU.scala 175:30]
  wire [7:0] _T_648 = ~(io_in_bits_Pctrl_adderRes_ori[58] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[47:40] :
    io_in_bits_DecodeIn_data_src2[47:40]; // @[PALU.scala 175:30]
  wire [7:0] _T_666 = ~(io_in_bits_Pctrl_adderRes_ori[68] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[55:48] :
    io_in_bits_DecodeIn_data_src2[55:48]; // @[PALU.scala 175:30]
  wire [7:0] _T_684 = ~(io_in_bits_Pctrl_adderRes_ori[78] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[63:56] :
    io_in_bits_DecodeIn_data_src2[63:56]; // @[PALU.scala 175:30]
  wire [63:0] _T_702 = {_T_684,_T_666,_T_648,_T_630,_T_612,_T_594,_T_576,_T_558}; // @[Cat.scala 30:58]
  wire  _T_705 = ~io_in_bits_DecodeIn_ctrl_funct3[1]; // @[PALU.scala 239:58]
  wire [63:0] _T_712 = ~(io_in_bits_Pctrl_adderRes_ori[64] ^ _T_705) ? io_in_bits_DecodeIn_data_src1 :
    io_in_bits_DecodeIn_data_src2; // @[PALU.scala 175:30]
  wire [31:0] _T_733 = ~(io_in_bits_Pctrl_adderRes_ori[32] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[31:0] :
    io_in_bits_DecodeIn_data_src2[31:0]; // @[PALU.scala 175:30]
  wire [31:0] _T_751 = ~(io_in_bits_Pctrl_adderRes_ori[66] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[63:32] :
    io_in_bits_DecodeIn_data_src2[63:32]; // @[PALU.scala 175:30]
  wire [63:0] _T_763 = {_T_751,_T_733}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_174 = io_in_bits_Pctrl_isMaxMin_32 ? _T_763 : 64'h0; // @[PALU.scala 240:28 241:19]
  wire [63:0] _GEN_175 = io_in_bits_Pctrl_isMaxMin_XLEN ? _T_712 : _GEN_174; // @[PALU.scala 238:30 239:19]
  wire [63:0] _GEN_176 = io_in_bits_Pctrl_isMaxMin_8 ? _T_702 : _GEN_175; // @[PALU.scala 236:27 237:19]
  wire [63:0] maxminRes = io_in_bits_Pctrl_isMaxMin_16 ? _T_548 : _GEN_176; // @[PALU.scala 234:22 235:19]
  wire [63:0] _T_766 = io_in_bits_DecodeIn_ctrl_fuOpType[0] ? io_in_bits_DecodeIn_data_src3 : 64'h0; // @[PALU.scala 247:22]
  wire [7:0] _T_770 = 8'hff ^ io_in_bits_Pctrl_adderRes[7:0]; // @[PALU.scala 247:128]
  wire [7:0] _T_772 = _T_770 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_774 = io_in_bits_Pctrl_adderRes_ori[8] ? _T_772 : io_in_bits_Pctrl_adderRes[7:0]; // @[PALU.scala 247:79]
  wire [7:0] _T_778 = 8'hff ^ io_in_bits_Pctrl_adderRes[15:8]; // @[PALU.scala 247:128]
  wire [7:0] _T_780 = _T_778 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_782 = io_in_bits_Pctrl_adderRes_ori[18] ? _T_780 : io_in_bits_Pctrl_adderRes[15:8]; // @[PALU.scala 247:79]
  wire [7:0] _T_786 = 8'hff ^ io_in_bits_Pctrl_adderRes[23:16]; // @[PALU.scala 247:128]
  wire [7:0] _T_788 = _T_786 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_790 = io_in_bits_Pctrl_adderRes_ori[28] ? _T_788 : io_in_bits_Pctrl_adderRes[23:16]; // @[PALU.scala 247:79]
  wire [7:0] _T_794 = 8'hff ^ io_in_bits_Pctrl_adderRes[31:24]; // @[PALU.scala 247:128]
  wire [7:0] _T_796 = _T_794 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_798 = io_in_bits_Pctrl_adderRes_ori[38] ? _T_796 : io_in_bits_Pctrl_adderRes[31:24]; // @[PALU.scala 247:79]
  wire [7:0] _T_802 = 8'hff ^ io_in_bits_Pctrl_adderRes[39:32]; // @[PALU.scala 247:128]
  wire [7:0] _T_804 = _T_802 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_806 = io_in_bits_Pctrl_adderRes_ori[48] ? _T_804 : io_in_bits_Pctrl_adderRes[39:32]; // @[PALU.scala 247:79]
  wire [7:0] _T_810 = 8'hff ^ io_in_bits_Pctrl_adderRes[47:40]; // @[PALU.scala 247:128]
  wire [7:0] _T_812 = _T_810 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_814 = io_in_bits_Pctrl_adderRes_ori[58] ? _T_812 : io_in_bits_Pctrl_adderRes[47:40]; // @[PALU.scala 247:79]
  wire [7:0] _T_818 = 8'hff ^ io_in_bits_Pctrl_adderRes[55:48]; // @[PALU.scala 247:128]
  wire [7:0] _T_820 = _T_818 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_822 = io_in_bits_Pctrl_adderRes_ori[68] ? _T_820 : io_in_bits_Pctrl_adderRes[55:48]; // @[PALU.scala 247:79]
  wire [7:0] _T_826 = 8'hff ^ io_in_bits_Pctrl_adderRes[63:56]; // @[PALU.scala 247:128]
  wire [7:0] _T_828 = _T_826 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_830 = io_in_bits_Pctrl_adderRes_ori[78] ? _T_828 : io_in_bits_Pctrl_adderRes[63:56]; // @[PALU.scala 247:79]
  wire [8:0] _T_831 = _T_774 + _T_782; // @[PALU.scala 247:188]
  wire [8:0] _GEN_648 = {{1'd0}, _T_790}; // @[PALU.scala 247:188]
  wire [9:0] _T_832 = _T_831 + _GEN_648; // @[PALU.scala 247:188]
  wire [9:0] _GEN_649 = {{2'd0}, _T_798}; // @[PALU.scala 247:188]
  wire [10:0] _T_833 = _T_832 + _GEN_649; // @[PALU.scala 247:188]
  wire [10:0] _GEN_650 = {{3'd0}, _T_806}; // @[PALU.scala 247:188]
  wire [11:0] _T_834 = _T_833 + _GEN_650; // @[PALU.scala 247:188]
  wire [11:0] _GEN_651 = {{4'd0}, _T_814}; // @[PALU.scala 247:188]
  wire [12:0] _T_835 = _T_834 + _GEN_651; // @[PALU.scala 247:188]
  wire [12:0] _GEN_652 = {{5'd0}, _T_822}; // @[PALU.scala 247:188]
  wire [13:0] _T_836 = _T_835 + _GEN_652; // @[PALU.scala 247:188]
  wire [13:0] _GEN_653 = {{6'd0}, _T_830}; // @[PALU.scala 247:188]
  wire [14:0] _T_837 = _T_836 + _GEN_653; // @[PALU.scala 247:188]
  wire [63:0] _GEN_654 = {{49'd0}, _T_837}; // @[PALU.scala 247:48]
  wire [63:0] _T_839 = _T_766 + _GEN_654; // @[PALU.scala 247:48]
  wire [63:0] pbsRes = io_in_bits_Pctrl_isPbs ? _T_839 : 64'h0; // @[PALU.scala 246:16 247:16]
  wire [4:0] _T_875 = 5'h1f ^ io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 367:52]
  wire [4:0] _T_877 = _T_875 + 5'h1; // @[PALU.scala 367:79]
  wire [4:0] _GEN_179 = _T_877 == 5'h10 ? 5'hf : _T_877; // @[PALU.scala 368:26 369:65 370:30]
  wire [4:0] _GEN_180 = io_in_bits_DecodeIn_data_src2[4] ? _GEN_179 : io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 366:47]
  wire [5:0] _T_884 = {io_in_bits_DecodeIn_data_src2[4],_GEN_180}; // @[Cat.scala 30:58]
  wire [3:0] _T_890 = 4'hf ^ io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 367:52]
  wire [3:0] _T_892 = _T_890 + 4'h1; // @[PALU.scala 367:79]
  wire [3:0] _GEN_182 = _T_892 == 4'h8 ? 4'h7 : _T_892; // @[PALU.scala 368:26 369:65 370:30]
  wire [3:0] _GEN_183 = io_in_bits_DecodeIn_data_src2[3] ? _GEN_182 : io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 366:47]
  wire [4:0] _T_899 = {io_in_bits_DecodeIn_data_src2[3],io_in_bits_DecodeIn_data_src2[3:0]}; // @[Cat.scala 30:58]
  wire [5:0] _T_900 = io_in_bits_Pctrl_isLR_16 ? _T_884 : {{1'd0}, _T_899}; // @[PALU.scala 500:22]
  wire [63:0] _WIRE_80 = {{58'd0}, _T_900};
  wire [4:0] _T_903 = io_in_bits_Pctrl_isLR_16 ? _WIRE_80[4:0] : {{1'd0}, _WIRE_80[3:0]}; // @[PALU.scala 501:27]
  wire  _T_907 = io_in_bits_Pctrl_isRs_16 | io_in_bits_Pctrl_isLR_16 & _WIRE_80[5]; // @[PALU.scala 503:70]
  wire [4:0] _T_911 = _T_903 - 5'h1; // @[PALU.scala 327:50]
  wire [4:0] _GEN_185 = io_in_bits_Pctrl_Round ? _T_911 : _T_903; // @[PALU.scala 327:{32,42}]
  wire [15:0] _T_912 = io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 329:42]
  wire [15:0] _T_914 = $signed(_T_912) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_915 = io_in_bits_DecodeIn_data_src1[15:0] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_186 = io_in_bits_Pctrl_Arithmetic ? _T_914 : _T_915; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_917 = {_GEN_186[15],_GEN_186}; // @[Cat.scala 30:58]
  wire [16:0] _T_918 = {1'h0,_GEN_186}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_187 = io_in_bits_Pctrl_Arithmetic ? _T_917 : _T_918; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_920 = _GEN_187 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_188 = io_in_bits_Pctrl_Round ? _T_920[16:1] : _GEN_186; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_931 = io_in_bits_DecodeIn_data_src1[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_932 = {_T_931,io_in_bits_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_2 = {{31'd0}, _T_932}; // @[PALU.scala 341:35]
  wire [62:0] _T_933 = _GEN_2 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_938 = 63'hffffffff ^ _T_933; // @[PALU.scala 345:80]
  wire [62:0] _GEN_189 = _T_933[31] ? _T_938 : _T_933; // @[PALU.scala 345:{53,59}]
  wire  _T_940 = _GEN_189[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_190 = _T_933[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_192 = _GEN_189[31:15] != 17'h0 ? _GEN_190 : _T_933[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_193 = io_in_bits_Pctrl_ShiftSigned & _T_940; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_194 = io_in_bits_Pctrl_ShiftSigned ? _GEN_192 : _T_933[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_195 = _T_907 ? _GEN_188 : _GEN_194; // @[PALU.scala 323:32]
  wire  _GEN_196 = _T_907 ? 1'h0 : _GEN_193; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_197 = _T_903 != 5'h0 ? _GEN_195 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_198 = _T_903 != 5'h0 & _GEN_196; // @[PALU.scala 322:31 317:45]
  wire [15:0] _T_966 = io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 329:42]
  wire [15:0] _T_968 = $signed(_T_966) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_969 = io_in_bits_DecodeIn_data_src1[31:16] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_200 = io_in_bits_Pctrl_Arithmetic ? _T_968 : _T_969; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_971 = {_GEN_200[15],_GEN_200}; // @[Cat.scala 30:58]
  wire [16:0] _T_972 = {1'h0,_GEN_200}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_201 = io_in_bits_Pctrl_Arithmetic ? _T_971 : _T_972; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_974 = _GEN_201 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_202 = io_in_bits_Pctrl_Round ? _T_974[16:1] : _GEN_200; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_985 = io_in_bits_DecodeIn_data_src1[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_986 = {_T_985,io_in_bits_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_4 = {{31'd0}, _T_986}; // @[PALU.scala 341:35]
  wire [62:0] _T_987 = _GEN_4 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_992 = 63'hffffffff ^ _T_987; // @[PALU.scala 345:80]
  wire [62:0] _GEN_203 = _T_987[31] ? _T_992 : _T_987; // @[PALU.scala 345:{53,59}]
  wire  _T_994 = _GEN_203[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_204 = _T_987[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_206 = _GEN_203[31:15] != 17'h0 ? _GEN_204 : _T_987[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_207 = io_in_bits_Pctrl_ShiftSigned & _T_994; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_208 = io_in_bits_Pctrl_ShiftSigned ? _GEN_206 : _T_987[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_209 = _T_907 ? _GEN_202 : _GEN_208; // @[PALU.scala 323:32]
  wire  _GEN_210 = _T_907 ? 1'h0 : _GEN_207; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_211 = _T_903 != 5'h0 ? _GEN_209 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_212 = _T_903 != 5'h0 & _GEN_210; // @[PALU.scala 322:31 317:45]
  wire [15:0] _T_1020 = io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 329:42]
  wire [15:0] _T_1022 = $signed(_T_1020) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_1023 = io_in_bits_DecodeIn_data_src1[47:32] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_214 = io_in_bits_Pctrl_Arithmetic ? _T_1022 : _T_1023; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_1025 = {_GEN_214[15],_GEN_214}; // @[Cat.scala 30:58]
  wire [16:0] _T_1026 = {1'h0,_GEN_214}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_215 = io_in_bits_Pctrl_Arithmetic ? _T_1025 : _T_1026; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_1028 = _GEN_215 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_216 = io_in_bits_Pctrl_Round ? _T_1028[16:1] : _GEN_214; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_1039 = io_in_bits_DecodeIn_data_src1[47] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1040 = {_T_1039,io_in_bits_DecodeIn_data_src1[47:32]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_6 = {{31'd0}, _T_1040}; // @[PALU.scala 341:35]
  wire [62:0] _T_1041 = _GEN_6 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_1046 = 63'hffffffff ^ _T_1041; // @[PALU.scala 345:80]
  wire [62:0] _GEN_217 = _T_1041[31] ? _T_1046 : _T_1041; // @[PALU.scala 345:{53,59}]
  wire  _T_1048 = _GEN_217[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_218 = _T_1041[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_220 = _GEN_217[31:15] != 17'h0 ? _GEN_218 : _T_1041[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_221 = io_in_bits_Pctrl_ShiftSigned & _T_1048; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_222 = io_in_bits_Pctrl_ShiftSigned ? _GEN_220 : _T_1041[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_223 = _T_907 ? _GEN_216 : _GEN_222; // @[PALU.scala 323:32]
  wire  _GEN_224 = _T_907 ? 1'h0 : _GEN_221; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_225 = _T_903 != 5'h0 ? _GEN_223 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_226 = _T_903 != 5'h0 & _GEN_224; // @[PALU.scala 322:31 317:45]
  wire [15:0] _T_1074 = io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 329:42]
  wire [15:0] _T_1076 = $signed(_T_1074) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_1077 = io_in_bits_DecodeIn_data_src1[63:48] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_228 = io_in_bits_Pctrl_Arithmetic ? _T_1076 : _T_1077; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_1079 = {_GEN_228[15],_GEN_228}; // @[Cat.scala 30:58]
  wire [16:0] _T_1080 = {1'h0,_GEN_228}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_229 = io_in_bits_Pctrl_Arithmetic ? _T_1079 : _T_1080; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_1082 = _GEN_229 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_230 = io_in_bits_Pctrl_Round ? _T_1082[16:1] : _GEN_228; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_1093 = io_in_bits_DecodeIn_data_src1[63] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1094 = {_T_1093,io_in_bits_DecodeIn_data_src1[63:48]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_9 = {{31'd0}, _T_1094}; // @[PALU.scala 341:35]
  wire [62:0] _T_1095 = _GEN_9 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_1100 = 63'hffffffff ^ _T_1095; // @[PALU.scala 345:80]
  wire [62:0] _GEN_231 = _T_1095[31] ? _T_1100 : _T_1095; // @[PALU.scala 345:{53,59}]
  wire  _T_1102 = _GEN_231[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_232 = _T_1095[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_234 = _GEN_231[31:15] != 17'h0 ? _GEN_232 : _T_1095[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_235 = io_in_bits_Pctrl_ShiftSigned & _T_1102; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_236 = io_in_bits_Pctrl_ShiftSigned ? _GEN_234 : _T_1095[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_237 = _T_907 ? _GEN_230 : _GEN_236; // @[PALU.scala 323:32]
  wire  _GEN_238 = _T_907 ? 1'h0 : _GEN_235; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_239 = _T_903 != 5'h0 ? _GEN_237 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_240 = _T_903 != 5'h0 & _GEN_238; // @[PALU.scala 322:31 317:45]
  wire  _T_1126 = _GEN_198 | _GEN_212 | _GEN_226 | _GEN_240; // @[PALU.scala 361:24]
  wire [64:0] _T_1130 = {_T_1126,_GEN_239,_GEN_225,_GEN_211,_GEN_197}; // @[Cat.scala 30:58]
  wire [4:0] _T_1150 = {io_in_bits_DecodeIn_data_src2[3],_GEN_183}; // @[Cat.scala 30:58]
  wire [3:0] _T_1165 = {io_in_bits_DecodeIn_data_src2[2],io_in_bits_DecodeIn_data_src2[2:0]}; // @[Cat.scala 30:58]
  wire [4:0] _T_1166 = io_in_bits_Pctrl_isLR_8 ? _T_1150 : {{1'd0}, _T_1165}; // @[PALU.scala 508:22]
  wire [63:0] _WIRE_120 = {{59'd0}, _T_1166};
  wire [3:0] _T_1169 = io_in_bits_Pctrl_isLR_8 ? _WIRE_120[3:0] : {{1'd0}, _WIRE_120[2:0]}; // @[PALU.scala 509:27]
  wire  _T_1173 = io_in_bits_Pctrl_isRs_8 | io_in_bits_Pctrl_isLR_8 & _WIRE_120[4]; // @[PALU.scala 511:68]
  wire [3:0] _T_1177 = _T_1169 - 4'h1; // @[PALU.scala 327:50]
  wire [3:0] _GEN_247 = io_in_bits_Pctrl_Round ? _T_1177 : _T_1169; // @[PALU.scala 327:{32,42}]
  wire [7:0] _T_1178 = io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 329:42]
  wire [7:0] _T_1180 = $signed(_T_1178) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1181 = io_in_bits_DecodeIn_data_src1[7:0] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_248 = io_in_bits_Pctrl_Arithmetic ? _T_1180 : _T_1181; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1183 = {_GEN_248[7],_GEN_248}; // @[Cat.scala 30:58]
  wire [8:0] _T_1184 = {1'h0,_GEN_248}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_249 = io_in_bits_Pctrl_Arithmetic ? _T_1183 : _T_1184; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1186 = _GEN_249 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_250 = io_in_bits_Pctrl_Round ? _T_1186[8:1] : _GEN_248; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1197 = io_in_bits_DecodeIn_data_src1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1198 = {_T_1197,io_in_bits_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_14 = {{15'd0}, _T_1198}; // @[PALU.scala 341:35]
  wire [30:0] _T_1199 = _GEN_14 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1204 = 31'hffff ^ _T_1199; // @[PALU.scala 345:80]
  wire [30:0] _GEN_251 = _T_1199[15] ? _T_1204 : _T_1199; // @[PALU.scala 345:{53,59}]
  wire  _T_1206 = _GEN_251[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_252 = _T_1199[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_254 = _GEN_251[15:7] != 9'h0 ? _GEN_252 : _T_1199[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_255 = io_in_bits_Pctrl_ShiftSigned & _T_1206; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_256 = io_in_bits_Pctrl_ShiftSigned ? _GEN_254 : _T_1199[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_257 = _T_1173 ? _GEN_250 : _GEN_256; // @[PALU.scala 323:32]
  wire  _GEN_258 = _T_1173 ? 1'h0 : _GEN_255; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_259 = _T_1169 != 4'h0 ? _GEN_257 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_260 = _T_1169 != 4'h0 & _GEN_258; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1232 = io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 329:42]
  wire [7:0] _T_1234 = $signed(_T_1232) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1235 = io_in_bits_DecodeIn_data_src1[15:8] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_262 = io_in_bits_Pctrl_Arithmetic ? _T_1234 : _T_1235; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1237 = {_GEN_262[7],_GEN_262}; // @[Cat.scala 30:58]
  wire [8:0] _T_1238 = {1'h0,_GEN_262}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_263 = io_in_bits_Pctrl_Arithmetic ? _T_1237 : _T_1238; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1240 = _GEN_263 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_264 = io_in_bits_Pctrl_Round ? _T_1240[8:1] : _GEN_262; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1251 = io_in_bits_DecodeIn_data_src1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1252 = {_T_1251,io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_16 = {{15'd0}, _T_1252}; // @[PALU.scala 341:35]
  wire [30:0] _T_1253 = _GEN_16 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1258 = 31'hffff ^ _T_1253; // @[PALU.scala 345:80]
  wire [30:0] _GEN_265 = _T_1253[15] ? _T_1258 : _T_1253; // @[PALU.scala 345:{53,59}]
  wire  _T_1260 = _GEN_265[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_266 = _T_1253[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_268 = _GEN_265[15:7] != 9'h0 ? _GEN_266 : _T_1253[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_269 = io_in_bits_Pctrl_ShiftSigned & _T_1260; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_270 = io_in_bits_Pctrl_ShiftSigned ? _GEN_268 : _T_1253[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_271 = _T_1173 ? _GEN_264 : _GEN_270; // @[PALU.scala 323:32]
  wire  _GEN_272 = _T_1173 ? 1'h0 : _GEN_269; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_273 = _T_1169 != 4'h0 ? _GEN_271 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_274 = _T_1169 != 4'h0 & _GEN_272; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1286 = io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 329:42]
  wire [7:0] _T_1288 = $signed(_T_1286) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1289 = io_in_bits_DecodeIn_data_src1[23:16] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_276 = io_in_bits_Pctrl_Arithmetic ? _T_1288 : _T_1289; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1291 = {_GEN_276[7],_GEN_276}; // @[Cat.scala 30:58]
  wire [8:0] _T_1292 = {1'h0,_GEN_276}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_277 = io_in_bits_Pctrl_Arithmetic ? _T_1291 : _T_1292; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1294 = _GEN_277 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_278 = io_in_bits_Pctrl_Round ? _T_1294[8:1] : _GEN_276; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1305 = io_in_bits_DecodeIn_data_src1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1306 = {_T_1305,io_in_bits_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_24 = {{15'd0}, _T_1306}; // @[PALU.scala 341:35]
  wire [30:0] _T_1307 = _GEN_24 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1312 = 31'hffff ^ _T_1307; // @[PALU.scala 345:80]
  wire [30:0] _GEN_279 = _T_1307[15] ? _T_1312 : _T_1307; // @[PALU.scala 345:{53,59}]
  wire  _T_1314 = _GEN_279[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_280 = _T_1307[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_282 = _GEN_279[15:7] != 9'h0 ? _GEN_280 : _T_1307[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_283 = io_in_bits_Pctrl_ShiftSigned & _T_1314; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_284 = io_in_bits_Pctrl_ShiftSigned ? _GEN_282 : _T_1307[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_285 = _T_1173 ? _GEN_278 : _GEN_284; // @[PALU.scala 323:32]
  wire  _GEN_286 = _T_1173 ? 1'h0 : _GEN_283; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_287 = _T_1169 != 4'h0 ? _GEN_285 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_288 = _T_1169 != 4'h0 & _GEN_286; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1340 = io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 329:42]
  wire [7:0] _T_1342 = $signed(_T_1340) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1343 = io_in_bits_DecodeIn_data_src1[31:24] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_290 = io_in_bits_Pctrl_Arithmetic ? _T_1342 : _T_1343; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1345 = {_GEN_290[7],_GEN_290}; // @[Cat.scala 30:58]
  wire [8:0] _T_1346 = {1'h0,_GEN_290}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_291 = io_in_bits_Pctrl_Arithmetic ? _T_1345 : _T_1346; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1348 = _GEN_291 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_292 = io_in_bits_Pctrl_Round ? _T_1348[8:1] : _GEN_290; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1359 = io_in_bits_DecodeIn_data_src1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1360 = {_T_1359,io_in_bits_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_26 = {{15'd0}, _T_1360}; // @[PALU.scala 341:35]
  wire [30:0] _T_1361 = _GEN_26 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1366 = 31'hffff ^ _T_1361; // @[PALU.scala 345:80]
  wire [30:0] _GEN_293 = _T_1361[15] ? _T_1366 : _T_1361; // @[PALU.scala 345:{53,59}]
  wire  _T_1368 = _GEN_293[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_294 = _T_1361[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_296 = _GEN_293[15:7] != 9'h0 ? _GEN_294 : _T_1361[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_297 = io_in_bits_Pctrl_ShiftSigned & _T_1368; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_298 = io_in_bits_Pctrl_ShiftSigned ? _GEN_296 : _T_1361[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_299 = _T_1173 ? _GEN_292 : _GEN_298; // @[PALU.scala 323:32]
  wire  _GEN_300 = _T_1173 ? 1'h0 : _GEN_297; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_301 = _T_1169 != 4'h0 ? _GEN_299 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_302 = _T_1169 != 4'h0 & _GEN_300; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1394 = io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 329:42]
  wire [7:0] _T_1396 = $signed(_T_1394) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1397 = io_in_bits_DecodeIn_data_src1[39:32] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_304 = io_in_bits_Pctrl_Arithmetic ? _T_1396 : _T_1397; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1399 = {_GEN_304[7],_GEN_304}; // @[Cat.scala 30:58]
  wire [8:0] _T_1400 = {1'h0,_GEN_304}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_305 = io_in_bits_Pctrl_Arithmetic ? _T_1399 : _T_1400; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1402 = _GEN_305 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_306 = io_in_bits_Pctrl_Round ? _T_1402[8:1] : _GEN_304; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1413 = io_in_bits_DecodeIn_data_src1[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1414 = {_T_1413,io_in_bits_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_34 = {{15'd0}, _T_1414}; // @[PALU.scala 341:35]
  wire [30:0] _T_1415 = _GEN_34 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1420 = 31'hffff ^ _T_1415; // @[PALU.scala 345:80]
  wire [30:0] _GEN_307 = _T_1415[15] ? _T_1420 : _T_1415; // @[PALU.scala 345:{53,59}]
  wire  _T_1422 = _GEN_307[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_308 = _T_1415[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_310 = _GEN_307[15:7] != 9'h0 ? _GEN_308 : _T_1415[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_311 = io_in_bits_Pctrl_ShiftSigned & _T_1422; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_312 = io_in_bits_Pctrl_ShiftSigned ? _GEN_310 : _T_1415[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_313 = _T_1173 ? _GEN_306 : _GEN_312; // @[PALU.scala 323:32]
  wire  _GEN_314 = _T_1173 ? 1'h0 : _GEN_311; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_315 = _T_1169 != 4'h0 ? _GEN_313 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_316 = _T_1169 != 4'h0 & _GEN_314; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1448 = io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 329:42]
  wire [7:0] _T_1450 = $signed(_T_1448) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1451 = io_in_bits_DecodeIn_data_src1[47:40] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_318 = io_in_bits_Pctrl_Arithmetic ? _T_1450 : _T_1451; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1453 = {_GEN_318[7],_GEN_318}; // @[Cat.scala 30:58]
  wire [8:0] _T_1454 = {1'h0,_GEN_318}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_319 = io_in_bits_Pctrl_Arithmetic ? _T_1453 : _T_1454; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1456 = _GEN_319 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_320 = io_in_bits_Pctrl_Round ? _T_1456[8:1] : _GEN_318; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1467 = io_in_bits_DecodeIn_data_src1[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1468 = {_T_1467,io_in_bits_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_36 = {{15'd0}, _T_1468}; // @[PALU.scala 341:35]
  wire [30:0] _T_1469 = _GEN_36 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1474 = 31'hffff ^ _T_1469; // @[PALU.scala 345:80]
  wire [30:0] _GEN_321 = _T_1469[15] ? _T_1474 : _T_1469; // @[PALU.scala 345:{53,59}]
  wire  _T_1476 = _GEN_321[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_322 = _T_1469[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_324 = _GEN_321[15:7] != 9'h0 ? _GEN_322 : _T_1469[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_325 = io_in_bits_Pctrl_ShiftSigned & _T_1476; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_326 = io_in_bits_Pctrl_ShiftSigned ? _GEN_324 : _T_1469[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_327 = _T_1173 ? _GEN_320 : _GEN_326; // @[PALU.scala 323:32]
  wire  _GEN_328 = _T_1173 ? 1'h0 : _GEN_325; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_329 = _T_1169 != 4'h0 ? _GEN_327 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_330 = _T_1169 != 4'h0 & _GEN_328; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1502 = io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 329:42]
  wire [7:0] _T_1504 = $signed(_T_1502) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1505 = io_in_bits_DecodeIn_data_src1[55:48] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_332 = io_in_bits_Pctrl_Arithmetic ? _T_1504 : _T_1505; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1507 = {_GEN_332[7],_GEN_332}; // @[Cat.scala 30:58]
  wire [8:0] _T_1508 = {1'h0,_GEN_332}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_333 = io_in_bits_Pctrl_Arithmetic ? _T_1507 : _T_1508; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1510 = _GEN_333 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_334 = io_in_bits_Pctrl_Round ? _T_1510[8:1] : _GEN_332; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1521 = io_in_bits_DecodeIn_data_src1[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1522 = {_T_1521,io_in_bits_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_45 = {{15'd0}, _T_1522}; // @[PALU.scala 341:35]
  wire [30:0] _T_1523 = _GEN_45 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1528 = 31'hffff ^ _T_1523; // @[PALU.scala 345:80]
  wire [30:0] _GEN_335 = _T_1523[15] ? _T_1528 : _T_1523; // @[PALU.scala 345:{53,59}]
  wire  _T_1530 = _GEN_335[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_336 = _T_1523[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_338 = _GEN_335[15:7] != 9'h0 ? _GEN_336 : _T_1523[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_339 = io_in_bits_Pctrl_ShiftSigned & _T_1530; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_340 = io_in_bits_Pctrl_ShiftSigned ? _GEN_338 : _T_1523[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_341 = _T_1173 ? _GEN_334 : _GEN_340; // @[PALU.scala 323:32]
  wire  _GEN_342 = _T_1173 ? 1'h0 : _GEN_339; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_343 = _T_1169 != 4'h0 ? _GEN_341 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_344 = _T_1169 != 4'h0 & _GEN_342; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1556 = io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 329:42]
  wire [7:0] _T_1558 = $signed(_T_1556) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1559 = io_in_bits_DecodeIn_data_src1[63:56] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_346 = io_in_bits_Pctrl_Arithmetic ? _T_1558 : _T_1559; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1561 = {_GEN_346[7],_GEN_346}; // @[Cat.scala 30:58]
  wire [8:0] _T_1562 = {1'h0,_GEN_346}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_347 = io_in_bits_Pctrl_Arithmetic ? _T_1561 : _T_1562; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1564 = _GEN_347 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_348 = io_in_bits_Pctrl_Round ? _T_1564[8:1] : _GEN_346; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1575 = io_in_bits_DecodeIn_data_src1[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1576 = {_T_1575,io_in_bits_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_47 = {{15'd0}, _T_1576}; // @[PALU.scala 341:35]
  wire [30:0] _T_1577 = _GEN_47 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1582 = 31'hffff ^ _T_1577; // @[PALU.scala 345:80]
  wire [30:0] _GEN_349 = _T_1577[15] ? _T_1582 : _T_1577; // @[PALU.scala 345:{53,59}]
  wire  _T_1584 = _GEN_349[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_350 = _T_1577[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_352 = _GEN_349[15:7] != 9'h0 ? _GEN_350 : _T_1577[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_353 = io_in_bits_Pctrl_ShiftSigned & _T_1584; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_354 = io_in_bits_Pctrl_ShiftSigned ? _GEN_352 : _T_1577[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_355 = _T_1173 ? _GEN_348 : _GEN_354; // @[PALU.scala 323:32]
  wire  _GEN_356 = _T_1173 ? 1'h0 : _GEN_353; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_357 = _T_1169 != 4'h0 ? _GEN_355 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_358 = _T_1169 != 4'h0 & _GEN_356; // @[PALU.scala 322:31 317:45]
  wire  _T_1612 = _GEN_260 | _GEN_274 | _GEN_288 | _GEN_302 | _GEN_316 | _GEN_330 | _GEN_344 | _GEN_358; // @[PALU.scala 361:24]
  wire [64:0] _T_1620 = {_T_1612,_GEN_357,_GEN_343,_GEN_329,_GEN_315,_GEN_301,_GEN_287,_GEN_273,_GEN_259}; // @[Cat.scala 30:58]
  wire  _T_1636 = io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isLR_32; // @[PALU.scala 517:32]
  wire [5:0] _T_1642 = 6'h3f ^ io_in_bits_DecodeIn_data_src2[5:0]; // @[PALU.scala 367:52]
  wire [5:0] _T_1644 = _T_1642 + 6'h1; // @[PALU.scala 367:79]
  wire [5:0] _GEN_359 = _T_1644 == 6'h20 ? 6'h1f : _T_1644; // @[PALU.scala 368:26 369:65 370:30]
  wire [5:0] _GEN_360 = io_in_bits_DecodeIn_data_src2[5] ? _GEN_359 : io_in_bits_DecodeIn_data_src2[5:0]; // @[PALU.scala 366:47]
  wire [6:0] _T_1651 = {io_in_bits_DecodeIn_data_src2[5],_GEN_360}; // @[Cat.scala 30:58]
  wire [5:0] _T_1666 = {io_in_bits_DecodeIn_data_src2[4],io_in_bits_DecodeIn_data_src2[4:0]}; // @[Cat.scala 30:58]
  wire [6:0] _T_1667 = io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isLR_32 ? _T_1651 : {{1'd0}, _T_1666}; // @[PALU.scala 517:22]
  wire [63:0] _WIRE_197 = {{57'd0}, _T_1667};
  wire [5:0] _T_1671 = _T_1636 ? _WIRE_197[5:0] : {{1'd0}, _WIRE_197[4:0]}; // @[PALU.scala 518:27]
  wire [63:0] _T_1675 = {32'h0,io_in_bits_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1676 = io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isLs_Q31 ? _T_1675 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 520:34]
  wire  _T_1681 = io_in_bits_Pctrl_isSRAIWU | io_in_bits_Pctrl_isRs_32 | (io_in_bits_Pctrl_isLR_32 |
    io_in_bits_Pctrl_isLR_Q31) & _WIRE_197[6]; // @[PALU.scala 520:130]
  wire [5:0] _T_1685 = _T_1671 - 6'h1; // @[PALU.scala 327:50]
  wire [5:0] _GEN_365 = io_in_bits_Pctrl_Round ? _T_1685 : _T_1671; // @[PALU.scala 327:{32,42}]
  wire [31:0] _T_1686 = _T_1676[31:0]; // @[PALU.scala 329:42]
  wire [31:0] _T_1688 = $signed(_T_1686) >>> _GEN_365; // @[PALU.scala 329:62]
  wire [31:0] _T_1689 = _T_1676[31:0] >> _GEN_365; // @[PALU.scala 331:41]
  wire [31:0] _GEN_366 = io_in_bits_Pctrl_Arithmetic ? _T_1688 : _T_1689; // @[PALU.scala 328:37 329:29 331:29]
  wire [32:0] _T_1691 = {_GEN_366[31],_GEN_366}; // @[Cat.scala 30:58]
  wire [32:0] _T_1692 = {1'h0,_GEN_366}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_367 = io_in_bits_Pctrl_Arithmetic ? _T_1691 : _T_1692; // @[PALU.scala 96:24 97:15 99:15]
  wire [32:0] _T_1694 = _GEN_367 + 33'h1; // @[PALU.scala 334:66]
  wire [31:0] _GEN_368 = io_in_bits_Pctrl_Round ? _T_1694[32:1] : _GEN_366; // @[PALU.scala 333:32 334:29 336:29]
  wire [31:0] _T_1705 = _T_1676[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1706 = {_T_1705,_T_1676[31:0]}; // @[Cat.scala 30:58]
  wire [126:0] _GEN_49 = {{63'd0}, _T_1706}; // @[PALU.scala 341:35]
  wire [126:0] _T_1707 = _GEN_49 << _T_1671; // @[PALU.scala 341:35]
  wire [126:0] _T_1712 = 127'hffffffffffffffff ^ _T_1707; // @[PALU.scala 345:80]
  wire [126:0] _GEN_369 = _T_1707[63] ? _T_1712 : _T_1707; // @[PALU.scala 345:{53,59}]
  wire  _T_1714 = _GEN_369[63:31] != 33'h0; // @[PALU.scala 346:54]
  wire [31:0] _GEN_370 = _T_1707[63] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 348:57 349:37 351:37]
  wire [31:0] _GEN_372 = _GEN_369[63:31] != 33'h0 ? _GEN_370 : _T_1707[31:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_373 = io_in_bits_Pctrl_ShiftSigned & _T_1714; // @[PALU.scala 343:38 317:45]
  wire [31:0] _GEN_374 = io_in_bits_Pctrl_ShiftSigned ? _GEN_372 : _T_1707[31:0]; // @[PALU.scala 342:25 343:38]
  wire [31:0] _GEN_375 = _T_1681 ? _GEN_368 : _GEN_374; // @[PALU.scala 323:32]
  wire  _GEN_376 = _T_1681 ? 1'h0 : _GEN_373; // @[PALU.scala 323:32 317:45]
  wire [31:0] _GEN_377 = _T_1671 != 6'h0 ? _GEN_375 : _T_1676[31:0]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_378 = _T_1671 != 6'h0 & _GEN_376; // @[PALU.scala 322:31 317:45]
  wire [31:0] _T_1740 = _T_1676[63:32]; // @[PALU.scala 329:42]
  wire [31:0] _T_1742 = $signed(_T_1740) >>> _GEN_365; // @[PALU.scala 329:62]
  wire [31:0] _T_1743 = _T_1676[63:32] >> _GEN_365; // @[PALU.scala 331:41]
  wire [31:0] _GEN_380 = io_in_bits_Pctrl_Arithmetic ? _T_1742 : _T_1743; // @[PALU.scala 328:37 329:29 331:29]
  wire [32:0] _T_1745 = {_GEN_380[31],_GEN_380}; // @[Cat.scala 30:58]
  wire [32:0] _T_1746 = {1'h0,_GEN_380}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_381 = io_in_bits_Pctrl_Arithmetic ? _T_1745 : _T_1746; // @[PALU.scala 96:24 97:15 99:15]
  wire [32:0] _T_1748 = _GEN_381 + 33'h1; // @[PALU.scala 334:66]
  wire [31:0] _GEN_382 = io_in_bits_Pctrl_Round ? _T_1748[32:1] : _GEN_380; // @[PALU.scala 333:32 334:29 336:29]
  wire [31:0] _T_1759 = _T_1676[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1760 = {_T_1759,_T_1676[63:32]}; // @[Cat.scala 30:58]
  wire [126:0] _GEN_52 = {{63'd0}, _T_1760}; // @[PALU.scala 341:35]
  wire [126:0] _T_1761 = _GEN_52 << _T_1671; // @[PALU.scala 341:35]
  wire [126:0] _T_1766 = 127'hffffffffffffffff ^ _T_1761; // @[PALU.scala 345:80]
  wire [126:0] _GEN_383 = _T_1761[63] ? _T_1766 : _T_1761; // @[PALU.scala 345:{53,59}]
  wire  _T_1768 = _GEN_383[63:31] != 33'h0; // @[PALU.scala 346:54]
  wire [31:0] _GEN_384 = _T_1761[63] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 348:57 349:37 351:37]
  wire [31:0] _GEN_386 = _GEN_383[63:31] != 33'h0 ? _GEN_384 : _T_1761[31:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_387 = io_in_bits_Pctrl_ShiftSigned & _T_1768; // @[PALU.scala 343:38 317:45]
  wire [31:0] _GEN_388 = io_in_bits_Pctrl_ShiftSigned ? _GEN_386 : _T_1761[31:0]; // @[PALU.scala 342:25 343:38]
  wire [31:0] _GEN_389 = _T_1681 ? _GEN_382 : _GEN_388; // @[PALU.scala 323:32]
  wire  _GEN_390 = _T_1681 ? 1'h0 : _GEN_387; // @[PALU.scala 323:32 317:45]
  wire [31:0] _GEN_391 = _T_1671 != 6'h0 ? _GEN_389 : _T_1676[63:32]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_392 = _T_1671 != 6'h0 & _GEN_390; // @[PALU.scala 322:31 317:45]
  wire  _T_1790 = _GEN_378 | _GEN_392; // @[PALU.scala 361:24]
  wire [64:0] _T_1792 = {_T_1790,_GEN_391,_GEN_377}; // @[Cat.scala 30:58]
  wire [31:0] _T_1798 = _T_1792[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1799 = {_T_1798,_T_1792[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1801 = io_in_bits_Pctrl_isLs_Q31 | io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isSRAIWU ? _T_1799 :
    _T_1792[63:0]; // @[PALU.scala 521:26]
  wire [6:0] _T_1827 = {io_in_bits_DecodeIn_data_src2[5],io_in_bits_DecodeIn_data_src2[5:0]}; // @[Cat.scala 30:58]
  wire [5:0] _T_1830 = io_in_bits_Pctrl_isRs_XLEN ? _T_1827[5:0] : {{1'd0}, _T_1827[4:0]}; // @[PALU.scala 526:27]
  wire [63:0] _T_1835 = {io_in_bits_DecodeIn_data_src1[31:0],io_in_bits_DecodeIn_data_src3[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1838 = {io_in_bits_DecodeIn_data_src3[31:0],io_in_bits_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1839 = _T_1827[5] ? _T_1835 : _T_1838; // @[PALU.scala 527:47]
  wire [63:0] _T_1840 = io_in_bits_Pctrl_isFSRW ? _T_1839 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 527:36]
  wire  _T_1841 = io_in_bits_Pctrl_isRs_XLEN & io_in_bits_Pctrl_Round; // @[PALU.scala 527:144]
  wire  _T_1843 = io_in_bits_Pctrl_isRs_XLEN & io_in_bits_Pctrl_Arithmetic; // @[PALU.scala 527:215]
  wire [5:0] _T_1847 = _T_1830 - 6'h1; // @[PALU.scala 327:50]
  wire [5:0] _GEN_396 = _T_1841 ? _T_1847 : _T_1830; // @[PALU.scala 327:{32,42}]
  wire [63:0] _T_1848 = io_in_bits_Pctrl_isFSRW ? _T_1839 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 329:42]
  wire [63:0] _T_1850 = $signed(_T_1848) >>> _GEN_396; // @[PALU.scala 329:62]
  wire [63:0] _T_1851 = _T_1840 >> _GEN_396; // @[PALU.scala 331:41]
  wire [63:0] _GEN_397 = _T_1843 ? _T_1850 : _T_1851; // @[PALU.scala 328:37 329:29 331:29]
  wire [64:0] _T_1853 = {_GEN_397[63],_GEN_397}; // @[Cat.scala 30:58]
  wire [64:0] _T_1854 = {1'h0,_GEN_397}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_398 = _T_1843 ? _T_1853 : _T_1854; // @[PALU.scala 96:24 97:15 99:15]
  wire [64:0] _T_1856 = _GEN_398 + 65'h1; // @[PALU.scala 334:66]
  wire [63:0] _GEN_399 = _T_1841 ? _T_1856[64:1] : _GEN_397; // @[PALU.scala 333:32 334:29 336:29]
  wire [63:0] _GEN_408 = _T_1830 != 6'h0 ? _GEN_399 : _T_1840; // @[PALU.scala 321:17 322:31]
  wire [64:0] _T_1898 = {1'h0,_GEN_408}; // @[Cat.scala 30:58]
  wire [31:0] _T_1903 = _T_1898[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1904 = {_T_1903,_T_1898[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1905 = io_in_bits_Pctrl_isRs_XLEN ? _T_1898[63:0] : _T_1904; // @[PALU.scala 528:26]
  wire [63:0] _GEN_410 = io_in_bits_Pctrl_isRs_XLEN | io_in_bits_Pctrl_isFSRW | io_in_bits_Pctrl_isWext ? _T_1905 :
    io_in_bits_DecodeIn_data_src1; // @[PALU.scala 524:44 528:20]
  wire  _GEN_411 = (io_in_bits_Pctrl_isRs_XLEN | io_in_bits_Pctrl_isFSRW | io_in_bits_Pctrl_isWext) & _T_1898[64]; // @[PALU.scala 524:44 529:20]
  wire [63:0] _GEN_412 = io_in_bits_Pctrl_isRs_32 | io_in_bits_Pctrl_isLs_32 | io_in_bits_Pctrl_isLR_32 |
    io_in_bits_Pctrl_isLs_Q31 | io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isSRAIWU ? _T_1801 : _GEN_410; // @[PALU.scala 515:77 521:20]
  wire  _GEN_413 = io_in_bits_Pctrl_isRs_32 | io_in_bits_Pctrl_isLs_32 | io_in_bits_Pctrl_isLR_32 |
    io_in_bits_Pctrl_isLs_Q31 | io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isSRAIWU ? _T_1792[64] : _GEN_411; // @[PALU.scala 515:77 522:20]
  wire [63:0] _GEN_414 = io_in_bits_Pctrl_isRs_8 | io_in_bits_Pctrl_isLs_8 | io_in_bits_Pctrl_isLR_8 ? _T_1620[63:0] :
    _GEN_412; // @[PALU.scala 506:40 512:20]
  wire  _GEN_415 = io_in_bits_Pctrl_isRs_8 | io_in_bits_Pctrl_isLs_8 | io_in_bits_Pctrl_isLR_8 ? _T_1620[64] : _GEN_413; // @[PALU.scala 506:40 513:20]
  wire [63:0] shifterRes = io_in_bits_Pctrl_isRs_16 | io_in_bits_Pctrl_isLs_16 | io_in_bits_Pctrl_isLR_16 ? _T_1130[63:0
    ] : _GEN_414; // @[PALU.scala 498:37 504:20]
  wire  shifterOV = io_in_bits_Pctrl_isRs_16 | io_in_bits_Pctrl_isLs_16 | io_in_bits_Pctrl_isLR_16 ? _T_1130[64] :
    _GEN_415; // @[PALU.scala 498:37 505:20]
  wire  _T_1909 = ~io_in_bits_DecodeIn_ctrl_func24; // @[PALU.scala 534:44]
  wire [15:0] _T_1914 = io_in_bits_DecodeIn_data_src1[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1916 = _T_1914 ^ io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_418 = _T_1909 ? _T_1916 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_1918 = _GEN_418 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire [30:0] _T_1920 = 31'hffff << io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 389:46]
  wire  _T_1921 = _T_1918 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_1925 = 16'hffff ^ _T_1920[15:0]; // @[PALU.scala 392:76]
  wire [15:0] _T_1926 = io_in_bits_DecodeIn_data_src1[15] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_1929 = ~_T_1909 & _T_1921; // @[PALU.scala 393:36]
  wire [15:0] _T_1933 = io_in_bits_DecodeIn_data_src1[15] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_420 = ~_T_1909 & _T_1921 ? _T_1933 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_421 = _T_1918 != 16'h0 & _T_1909 | _T_1929; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_422 = _T_1918 != 16'h0 & _T_1909 ? _T_1926 : _GEN_420; // @[PALU.scala 390:44 392:21]
  wire [15:0] _T_1945 = io_in_bits_DecodeIn_data_src1[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1947 = _T_1945 ^ io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_423 = _T_1909 ? _T_1947 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_1949 = _GEN_423 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire  _T_1952 = _T_1949 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_1957 = io_in_bits_DecodeIn_data_src1[31] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_1960 = ~_T_1909 & _T_1952; // @[PALU.scala 393:36]
  wire [15:0] _T_1964 = io_in_bits_DecodeIn_data_src1[31] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_425 = ~_T_1909 & _T_1952 ? _T_1964 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_426 = _T_1949 != 16'h0 & _T_1909 | _T_1960; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_427 = _T_1949 != 16'h0 & _T_1909 ? _T_1957 : _GEN_425; // @[PALU.scala 390:44 392:21]
  wire [15:0] _T_1976 = io_in_bits_DecodeIn_data_src1[47] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1978 = _T_1976 ^ io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_428 = _T_1909 ? _T_1978 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_1980 = _GEN_428 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire  _T_1983 = _T_1980 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_1988 = io_in_bits_DecodeIn_data_src1[47] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_1991 = ~_T_1909 & _T_1983; // @[PALU.scala 393:36]
  wire [15:0] _T_1995 = io_in_bits_DecodeIn_data_src1[47] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_430 = ~_T_1909 & _T_1983 ? _T_1995 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_431 = _T_1980 != 16'h0 & _T_1909 | _T_1991; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_432 = _T_1980 != 16'h0 & _T_1909 ? _T_1988 : _GEN_430; // @[PALU.scala 390:44 392:21]
  wire [15:0] _T_2007 = io_in_bits_DecodeIn_data_src1[63] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2009 = _T_2007 ^ io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_433 = _T_1909 ? _T_2009 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_2011 = _GEN_433 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire  _T_2014 = _T_2011 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_2019 = io_in_bits_DecodeIn_data_src1[63] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_2022 = ~_T_1909 & _T_2014; // @[PALU.scala 393:36]
  wire [15:0] _T_2026 = io_in_bits_DecodeIn_data_src1[63] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_435 = ~_T_1909 & _T_2014 ? _T_2026 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_436 = _T_2011 != 16'h0 & _T_1909 | _T_2022; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_437 = _T_2011 != 16'h0 & _T_1909 ? _T_2019 : _GEN_435; // @[PALU.scala 390:44 392:21]
  wire  _T_2036 = _GEN_421 | _GEN_426 | _GEN_431 | _GEN_436; // @[PALU.scala 400:24]
  wire [64:0] _T_2040 = {_T_2036,_GEN_437,_GEN_432,_GEN_427,_GEN_422}; // @[Cat.scala 30:58]
  wire [7:0] _T_2049 = io_in_bits_DecodeIn_data_src1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2051 = _T_2049 ^ io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_438 = _T_1909 ? _T_2051 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2053 = _GEN_438 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire [14:0] _T_2055 = 15'hff << io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 389:46]
  wire  _T_2056 = _T_2053 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2060 = 8'hff ^ _T_2055[7:0]; // @[PALU.scala 392:76]
  wire [7:0] _T_2061 = io_in_bits_DecodeIn_data_src1[7] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2064 = ~_T_1909 & _T_2056; // @[PALU.scala 393:36]
  wire [7:0] _T_2068 = io_in_bits_DecodeIn_data_src1[7] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_440 = ~_T_1909 & _T_2056 ? _T_2068 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_441 = _T_2053 != 8'h0 & _T_1909 | _T_2064; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_442 = _T_2053 != 8'h0 & _T_1909 ? _T_2061 : _GEN_440; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2080 = io_in_bits_DecodeIn_data_src1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2082 = _T_2080 ^ io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_443 = _T_1909 ? _T_2082 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2084 = _GEN_443 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2087 = _T_2084 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2092 = io_in_bits_DecodeIn_data_src1[15] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2095 = ~_T_1909 & _T_2087; // @[PALU.scala 393:36]
  wire [7:0] _T_2099 = io_in_bits_DecodeIn_data_src1[15] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_445 = ~_T_1909 & _T_2087 ? _T_2099 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_446 = _T_2084 != 8'h0 & _T_1909 | _T_2095; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_447 = _T_2084 != 8'h0 & _T_1909 ? _T_2092 : _GEN_445; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2111 = io_in_bits_DecodeIn_data_src1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2113 = _T_2111 ^ io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_448 = _T_1909 ? _T_2113 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2115 = _GEN_448 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2118 = _T_2115 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2123 = io_in_bits_DecodeIn_data_src1[23] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2126 = ~_T_1909 & _T_2118; // @[PALU.scala 393:36]
  wire [7:0] _T_2130 = io_in_bits_DecodeIn_data_src1[23] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_450 = ~_T_1909 & _T_2118 ? _T_2130 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_451 = _T_2115 != 8'h0 & _T_1909 | _T_2126; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_452 = _T_2115 != 8'h0 & _T_1909 ? _T_2123 : _GEN_450; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2142 = io_in_bits_DecodeIn_data_src1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2144 = _T_2142 ^ io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_453 = _T_1909 ? _T_2144 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2146 = _GEN_453 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2149 = _T_2146 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2154 = io_in_bits_DecodeIn_data_src1[31] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2157 = ~_T_1909 & _T_2149; // @[PALU.scala 393:36]
  wire [7:0] _T_2161 = io_in_bits_DecodeIn_data_src1[31] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_455 = ~_T_1909 & _T_2149 ? _T_2161 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_456 = _T_2146 != 8'h0 & _T_1909 | _T_2157; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_457 = _T_2146 != 8'h0 & _T_1909 ? _T_2154 : _GEN_455; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2173 = io_in_bits_DecodeIn_data_src1[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2175 = _T_2173 ^ io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_458 = _T_1909 ? _T_2175 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2177 = _GEN_458 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2180 = _T_2177 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2185 = io_in_bits_DecodeIn_data_src1[39] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2188 = ~_T_1909 & _T_2180; // @[PALU.scala 393:36]
  wire [7:0] _T_2192 = io_in_bits_DecodeIn_data_src1[39] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_460 = ~_T_1909 & _T_2180 ? _T_2192 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_461 = _T_2177 != 8'h0 & _T_1909 | _T_2188; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_462 = _T_2177 != 8'h0 & _T_1909 ? _T_2185 : _GEN_460; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2204 = io_in_bits_DecodeIn_data_src1[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2206 = _T_2204 ^ io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_463 = _T_1909 ? _T_2206 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2208 = _GEN_463 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2211 = _T_2208 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2216 = io_in_bits_DecodeIn_data_src1[47] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2219 = ~_T_1909 & _T_2211; // @[PALU.scala 393:36]
  wire [7:0] _T_2223 = io_in_bits_DecodeIn_data_src1[47] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_465 = ~_T_1909 & _T_2211 ? _T_2223 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_466 = _T_2208 != 8'h0 & _T_1909 | _T_2219; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_467 = _T_2208 != 8'h0 & _T_1909 ? _T_2216 : _GEN_465; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2235 = io_in_bits_DecodeIn_data_src1[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2237 = _T_2235 ^ io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_468 = _T_1909 ? _T_2237 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2239 = _GEN_468 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2242 = _T_2239 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2247 = io_in_bits_DecodeIn_data_src1[55] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2250 = ~_T_1909 & _T_2242; // @[PALU.scala 393:36]
  wire [7:0] _T_2254 = io_in_bits_DecodeIn_data_src1[55] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_470 = ~_T_1909 & _T_2242 ? _T_2254 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_471 = _T_2239 != 8'h0 & _T_1909 | _T_2250; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_472 = _T_2239 != 8'h0 & _T_1909 ? _T_2247 : _GEN_470; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2266 = io_in_bits_DecodeIn_data_src1[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2268 = _T_2266 ^ io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_473 = _T_1909 ? _T_2268 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2270 = _GEN_473 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2273 = _T_2270 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2278 = io_in_bits_DecodeIn_data_src1[63] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2281 = ~_T_1909 & _T_2273; // @[PALU.scala 393:36]
  wire [7:0] _T_2285 = io_in_bits_DecodeIn_data_src1[63] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_475 = ~_T_1909 & _T_2273 ? _T_2285 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_476 = _T_2270 != 8'h0 & _T_1909 | _T_2281; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_477 = _T_2270 != 8'h0 & _T_1909 ? _T_2278 : _GEN_475; // @[PALU.scala 390:44 392:21]
  wire  _T_2299 = _GEN_441 | _GEN_446 | _GEN_451 | _GEN_456 | _GEN_461 | _GEN_466 | _GEN_471 | _GEN_476; // @[PALU.scala 400:24]
  wire [64:0] _T_2307 = {_T_2299,_GEN_477,_GEN_472,_GEN_467,_GEN_462,_GEN_457,_GEN_452,_GEN_447,_GEN_442}; // @[Cat.scala 30:58]
  wire [31:0] _T_2317 = io_in_bits_DecodeIn_data_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2319 = _T_2317 ^ io_in_bits_DecodeIn_data_src1[31:0]; // @[PALU.scala 384:58]
  wire [31:0] _GEN_478 = _T_15 ? _T_2319 : io_in_bits_DecodeIn_data_src1[31:0]; // @[PALU.scala 383:29 384:22 386:22]
  wire [31:0] _T_2321 = _GEN_478 >> io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 388:28]
  wire [62:0] _T_2323 = 63'hffffffff << io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 389:46]
  wire  _T_2324 = _T_2321 != 32'h0; // @[PALU.scala 390:22]
  wire [31:0] _T_2328 = 32'hffffffff ^ _T_2323[31:0]; // @[PALU.scala 392:76]
  wire [31:0] _T_2329 = io_in_bits_DecodeIn_data_src1[31] ? _T_2323[31:0] : _T_2328; // @[PALU.scala 392:27]
  wire  _T_2332 = ~_T_15 & _T_2324; // @[PALU.scala 393:36]
  wire [31:0] _T_2336 = io_in_bits_DecodeIn_data_src1[31] ? 32'h0 : _T_2328; // @[PALU.scala 395:27]
  wire [31:0] _GEN_480 = ~_T_15 & _T_2324 ? _T_2336 : io_in_bits_DecodeIn_data_src1[31:0]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_481 = _T_2321 != 32'h0 & _T_15 | _T_2332; // @[PALU.scala 390:44 391:23]
  wire [31:0] _GEN_482 = _T_2321 != 32'h0 & _T_15 ? _T_2329 : _GEN_480; // @[PALU.scala 390:44 392:21]
  wire [31:0] _T_2348 = io_in_bits_DecodeIn_data_src1[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2350 = _T_2348 ^ io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 384:58]
  wire [31:0] _GEN_483 = _T_15 ? _T_2350 : io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 383:29 384:22 386:22]
  wire [31:0] _T_2352 = _GEN_483 >> io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 388:28]
  wire  _T_2355 = _T_2352 != 32'h0; // @[PALU.scala 390:22]
  wire [31:0] _T_2360 = io_in_bits_DecodeIn_data_src1[63] ? _T_2323[31:0] : _T_2328; // @[PALU.scala 392:27]
  wire  _T_2363 = ~_T_15 & _T_2355; // @[PALU.scala 393:36]
  wire [31:0] _T_2367 = io_in_bits_DecodeIn_data_src1[63] ? 32'h0 : _T_2328; // @[PALU.scala 395:27]
  wire [31:0] _GEN_485 = ~_T_15 & _T_2355 ? _T_2367 : io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_486 = _T_2352 != 32'h0 & _T_15 | _T_2363; // @[PALU.scala 390:44 391:23]
  wire [31:0] _GEN_487 = _T_2352 != 32'h0 & _T_15 ? _T_2360 : _GEN_485; // @[PALU.scala 390:44 392:21]
  wire  _T_2375 = _GEN_481 | _GEN_486; // @[PALU.scala 400:24]
  wire [64:0] _T_2377 = {_T_2375,_GEN_487,_GEN_482}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_488 = io_in_bits_Pctrl_isclip_32 ? _T_2377[63:0] : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 541:26 543:17]
  wire  _GEN_489 = io_in_bits_Pctrl_isclip_32 & _T_2377[64]; // @[PALU.scala 541:26 544:17]
  wire [63:0] _GEN_490 = io_in_bits_Pctrl_isClip_8 ? _T_2307[63:0] : _GEN_488; // @[PALU.scala 537:25 539:17]
  wire  _GEN_491 = io_in_bits_Pctrl_isClip_8 ? _T_2307[64] : _GEN_489; // @[PALU.scala 537:25 540:17]
  wire [63:0] clipRes = io_in_bits_Pctrl_isClip_16 ? _T_2040[63:0] : _GEN_490; // @[PALU.scala 533:20 535:17]
  wire  clipOV = io_in_bits_Pctrl_isClip_16 ? _T_2040[64] : _GEN_491; // @[PALU.scala 533:20 536:17]
  wire  _T_2384 = io_in_bits_DecodeIn_data_src1[15:0] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2390 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 413:42]
  wire [15:0] _T_2392 = _T_2390 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_494 = io_in_bits_DecodeIn_data_src1[15] ? _T_2392 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_496 = io_in_bits_DecodeIn_data_src1[15:0] == 16'h8000 ? 16'h7fff : _GEN_494; // @[PALU.scala 409:53 411:23]
  wire  _T_2397 = io_in_bits_DecodeIn_data_src1[31:16] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2403 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 413:42]
  wire [15:0] _T_2405 = _T_2403 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_497 = io_in_bits_DecodeIn_data_src1[31] ? _T_2405 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_499 = io_in_bits_DecodeIn_data_src1[31:16] == 16'h8000 ? 16'h7fff : _GEN_497; // @[PALU.scala 409:53 411:23]
  wire  _T_2410 = io_in_bits_DecodeIn_data_src1[47:32] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2416 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 413:42]
  wire [15:0] _T_2418 = _T_2416 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_500 = io_in_bits_DecodeIn_data_src1[47] ? _T_2418 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_502 = io_in_bits_DecodeIn_data_src1[47:32] == 16'h8000 ? 16'h7fff : _GEN_500; // @[PALU.scala 409:53 411:23]
  wire  _T_2423 = io_in_bits_DecodeIn_data_src1[63:48] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2429 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 413:42]
  wire [15:0] _T_2431 = _T_2429 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_503 = io_in_bits_DecodeIn_data_src1[63] ? _T_2431 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_505 = io_in_bits_DecodeIn_data_src1[63:48] == 16'h8000 ? 16'h7fff : _GEN_503; // @[PALU.scala 409:53 411:23]
  wire  _T_2434 = _T_2384 | _T_2397 | _T_2410 | _T_2423; // @[PALU.scala 417:24]
  wire [64:0] _T_2438 = {_T_2434,_GEN_505,_GEN_502,_GEN_499,_GEN_496}; // @[Cat.scala 30:58]
  wire  _T_2445 = io_in_bits_DecodeIn_data_src1[7:0] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2451 = 8'hff ^ io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 413:42]
  wire [7:0] _T_2453 = _T_2451 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_506 = io_in_bits_DecodeIn_data_src1[7] ? _T_2453 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_508 = io_in_bits_DecodeIn_data_src1[7:0] == 8'h80 ? 8'h7f : _GEN_506; // @[PALU.scala 409:53 411:23]
  wire  _T_2458 = io_in_bits_DecodeIn_data_src1[15:8] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2464 = 8'hff ^ io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 413:42]
  wire [7:0] _T_2466 = _T_2464 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_509 = io_in_bits_DecodeIn_data_src1[15] ? _T_2466 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_511 = io_in_bits_DecodeIn_data_src1[15:8] == 8'h80 ? 8'h7f : _GEN_509; // @[PALU.scala 409:53 411:23]
  wire  _T_2471 = io_in_bits_DecodeIn_data_src1[23:16] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2477 = 8'hff ^ io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 413:42]
  wire [7:0] _T_2479 = _T_2477 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_512 = io_in_bits_DecodeIn_data_src1[23] ? _T_2479 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_514 = io_in_bits_DecodeIn_data_src1[23:16] == 8'h80 ? 8'h7f : _GEN_512; // @[PALU.scala 409:53 411:23]
  wire  _T_2484 = io_in_bits_DecodeIn_data_src1[31:24] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2490 = 8'hff ^ io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 413:42]
  wire [7:0] _T_2492 = _T_2490 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_515 = io_in_bits_DecodeIn_data_src1[31] ? _T_2492 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_517 = io_in_bits_DecodeIn_data_src1[31:24] == 8'h80 ? 8'h7f : _GEN_515; // @[PALU.scala 409:53 411:23]
  wire  _T_2497 = io_in_bits_DecodeIn_data_src1[39:32] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2503 = 8'hff ^ io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 413:42]
  wire [7:0] _T_2505 = _T_2503 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_518 = io_in_bits_DecodeIn_data_src1[39] ? _T_2505 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_520 = io_in_bits_DecodeIn_data_src1[39:32] == 8'h80 ? 8'h7f : _GEN_518; // @[PALU.scala 409:53 411:23]
  wire  _T_2510 = io_in_bits_DecodeIn_data_src1[47:40] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2516 = 8'hff ^ io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 413:42]
  wire [7:0] _T_2518 = _T_2516 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_521 = io_in_bits_DecodeIn_data_src1[47] ? _T_2518 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_523 = io_in_bits_DecodeIn_data_src1[47:40] == 8'h80 ? 8'h7f : _GEN_521; // @[PALU.scala 409:53 411:23]
  wire  _T_2523 = io_in_bits_DecodeIn_data_src1[55:48] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2529 = 8'hff ^ io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 413:42]
  wire [7:0] _T_2531 = _T_2529 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_524 = io_in_bits_DecodeIn_data_src1[55] ? _T_2531 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_526 = io_in_bits_DecodeIn_data_src1[55:48] == 8'h80 ? 8'h7f : _GEN_524; // @[PALU.scala 409:53 411:23]
  wire  _T_2536 = io_in_bits_DecodeIn_data_src1[63:56] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2542 = 8'hff ^ io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 413:42]
  wire [7:0] _T_2544 = _T_2542 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_527 = io_in_bits_DecodeIn_data_src1[63] ? _T_2544 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_529 = io_in_bits_DecodeIn_data_src1[63:56] == 8'h80 ? 8'h7f : _GEN_527; // @[PALU.scala 409:53 411:23]
  wire  _T_2551 = _T_2445 | _T_2458 | _T_2471 | _T_2484 | _T_2497 | _T_2510 | _T_2523 | _T_2536; // @[PALU.scala 417:24]
  wire [64:0] _T_2559 = {_T_2551,_GEN_529,_GEN_526,_GEN_523,_GEN_520,_GEN_517,_GEN_514,_GEN_511,_GEN_508}; // @[Cat.scala 30:58]
  wire [63:0] _T_2565 = io_in_bits_Pctrl_isSat_W ? _T_1675 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 558:35]
  wire  _T_2570 = _T_2565[31:0] == 32'h80000000; // @[PALU.scala 409:22]
  wire [31:0] _T_2576 = 32'hffffffff ^ _T_2565[31:0]; // @[PALU.scala 413:42]
  wire [31:0] _T_2578 = _T_2576 + 32'h1; // @[PALU.scala 413:48]
  wire [31:0] _GEN_530 = _T_2565[31] ? _T_2578 : _T_2565[31:0]; // @[PALU.scala 412:44 413:23]
  wire [31:0] _GEN_532 = _T_2565[31:0] == 32'h80000000 ? 32'h7fffffff : _GEN_530; // @[PALU.scala 409:53 411:23]
  wire  _T_2583 = _T_2565[63:32] == 32'h80000000; // @[PALU.scala 409:22]
  wire [31:0] _T_2589 = 32'hffffffff ^ _T_2565[63:32]; // @[PALU.scala 413:42]
  wire [31:0] _T_2591 = _T_2589 + 32'h1; // @[PALU.scala 413:48]
  wire [31:0] _GEN_533 = _T_2565[63] ? _T_2591 : _T_2565[63:32]; // @[PALU.scala 412:44 413:23]
  wire [31:0] _GEN_535 = _T_2565[63:32] == 32'h80000000 ? 32'h7fffffff : _GEN_533; // @[PALU.scala 409:53 411:23]
  wire  _T_2592 = _T_2570 | _T_2583; // @[PALU.scala 417:24]
  wire [64:0] _T_2594 = {_T_2592,_GEN_535,_GEN_532}; // @[Cat.scala 30:58]
  wire [31:0] _T_2598 = _T_2594[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2599 = {_T_2598,_T_2594[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2601 = io_in_bits_Pctrl_isSat_W ? _T_2599 : _T_2594[63:0]; // @[PALU.scala 559:22]
  wire [63:0] _GEN_536 = io_in_bits_Pctrl_isSat_32 | io_in_bits_Pctrl_isSat_W ? _T_2601 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 557:35 559:16]
  wire  _GEN_537 = (io_in_bits_Pctrl_isSat_32 | io_in_bits_Pctrl_isSat_W) & _T_2594[64]; // @[PALU.scala 557:35 560:16]
  wire [63:0] _GEN_538 = io_in_bits_Pctrl_isSat_8 ? _T_2559[63:0] : _GEN_536; // @[PALU.scala 553:24 555:16]
  wire  _GEN_539 = io_in_bits_Pctrl_isSat_8 ? _T_2559[64] : _GEN_537; // @[PALU.scala 553:24 556:16]
  wire [63:0] satRes = io_in_bits_Pctrl_isSat_16 ? _T_2438[63:0] : _GEN_538; // @[PALU.scala 549:19 551:16]
  wire  satOV = io_in_bits_Pctrl_isSat_16 ? _T_2438[64] : _GEN_539; // @[PALU.scala 549:19 552:16]
  wire [4:0] _T_2604 = io_in_bits_DecodeIn_data_src2[4:0] & 5'h1b; // @[PALU.scala 566:45]
  wire  _T_2607 = ~io_in_bits_DecodeIn_data_src2[2]; // @[PALU.scala 566:57]
  wire [7:0] _T_2616 = io_in_bits_DecodeIn_data_src1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2617 = {_T_2616,io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2618 = {8'h0,io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_542 = _T_2607 ? _T_2617 : _T_2618; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2626 = io_in_bits_DecodeIn_data_src1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2627 = {_T_2626,io_in_bits_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2628 = {8'h0,io_in_bits_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_543 = _T_2607 ? _T_2627 : _T_2628; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2635 = io_in_bits_DecodeIn_data_src1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2636 = {_T_2635,io_in_bits_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2637 = {8'h0,io_in_bits_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_544 = _T_2607 ? _T_2636 : _T_2637; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2638 = _T_2604 == 5'h9 ? _GEN_543 : _GEN_544; // @[PALU.scala 464:107]
  wire [15:0] _T_2639 = _T_2604 == 5'h8 ? _GEN_542 : _T_2638; // @[PALU.scala 464:26]
  wire [7:0] _T_2666 = io_in_bits_DecodeIn_data_src1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2667 = {_T_2666,io_in_bits_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2668 = {8'h0,io_in_bits_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_547 = _T_2607 ? _T_2667 : _T_2668; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2669 = _T_2604 == 5'hb ? _GEN_542 : _GEN_547; // @[PALU.scala 465:107]
  wire [15:0] _T_2670 = _T_2604 == 5'h13 ? _GEN_543 : _T_2669; // @[PALU.scala 465:26]
  wire [7:0] _T_2680 = io_in_bits_DecodeIn_data_src1[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2681 = {_T_2680,io_in_bits_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2682 = {8'h0,io_in_bits_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_548 = _T_2607 ? _T_2681 : _T_2682; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2690 = io_in_bits_DecodeIn_data_src1[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2691 = {_T_2690,io_in_bits_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2692 = {8'h0,io_in_bits_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_549 = _T_2607 ? _T_2691 : _T_2692; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2699 = io_in_bits_DecodeIn_data_src1[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2700 = {_T_2699,io_in_bits_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2701 = {8'h0,io_in_bits_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_550 = _T_2607 ? _T_2700 : _T_2701; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2702 = _T_2604 == 5'h9 ? _GEN_549 : _GEN_550; // @[PALU.scala 464:107]
  wire [15:0] _T_2703 = _T_2604 == 5'h8 ? _GEN_548 : _T_2702; // @[PALU.scala 464:26]
  wire [7:0] _T_2730 = io_in_bits_DecodeIn_data_src1[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2731 = {_T_2730,io_in_bits_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2732 = {8'h0,io_in_bits_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_553 = _T_2607 ? _T_2731 : _T_2732; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2733 = _T_2604 == 5'hb ? _GEN_548 : _GEN_553; // @[PALU.scala 465:107]
  wire [15:0] _T_2734 = _T_2604 == 5'h13 ? _GEN_549 : _T_2733; // @[PALU.scala 465:26]
  wire [63:0] _T_2736 = {_T_2703,_T_2734,_T_2639,_T_2670}; // @[Cat.scala 30:58]
  wire [63:0] unpackRes = io_in_bits_Pctrl_isUnpack ? _T_2736 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 565:19 566:19]
  wire  _T_2740 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[15]; // @[PALU.scala 423:29]
  wire  _T_2742 = io_in_bits_DecodeIn_data_src1[0] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2744 = io_in_bits_DecodeIn_data_src1[1] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2746 = io_in_bits_DecodeIn_data_src1[2] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2748 = io_in_bits_DecodeIn_data_src1[3] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2750 = io_in_bits_DecodeIn_data_src1[4] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2752 = io_in_bits_DecodeIn_data_src1[5] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2754 = io_in_bits_DecodeIn_data_src1[6] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2756 = io_in_bits_DecodeIn_data_src1[7] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2758 = io_in_bits_DecodeIn_data_src1[8] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2760 = io_in_bits_DecodeIn_data_src1[9] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2762 = io_in_bits_DecodeIn_data_src1[10] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2764 = io_in_bits_DecodeIn_data_src1[11] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2766 = io_in_bits_DecodeIn_data_src1[12] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2768 = io_in_bits_DecodeIn_data_src1[13] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2770 = io_in_bits_DecodeIn_data_src1[14] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2772 = io_in_bits_DecodeIn_data_src1[15] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2774 = _T_2770 & _T_2772; // @[PALU.scala 427:113]
  wire  _T_2776 = _T_2768 & (_T_2770 & _T_2772); // @[PALU.scala 427:113]
  wire  _T_2778 = _T_2766 & (_T_2768 & (_T_2770 & _T_2772)); // @[PALU.scala 427:113]
  wire  _T_2780 = _T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))); // @[PALU.scala 427:113]
  wire  _T_2782 = _T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))); // @[PALU.scala 427:113]
  wire  _T_2784 = _T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))))); // @[PALU.scala 427:113]
  wire  _T_2786 = _T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))))); // @[PALU.scala 427:113]
  wire  _T_2788 = _T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))))))); // @[PALU.scala 427:113]
  wire  _T_2790 = _T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 &
    _T_2772)))))))); // @[PALU.scala 427:113]
  wire  _T_2792 = _T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (
    _T_2770 & _T_2772))))))))); // @[PALU.scala 427:113]
  wire  _T_2794 = _T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (
    _T_2768 & (_T_2770 & _T_2772)))))))))); // @[PALU.scala 427:113]
  wire  _T_2796 = _T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (
    _T_2766 & (_T_2768 & (_T_2770 & _T_2772))))))))))); // @[PALU.scala 427:113]
  wire  _T_2798 = _T_2746 & (_T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (
    _T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))))))))))); // @[PALU.scala 427:113]
  wire  _T_2800 = _T_2744 & (_T_2746 & (_T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (
    _T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))))))))))))); // @[PALU.scala 427:113]
  wire  _T_2802 = _T_2742 & (_T_2744 & (_T_2746 & (_T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (
    _T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_2803 = _T_2772 + _T_2774; // @[PALU.scala 428:38]
  wire [1:0] _GEN_655 = {{1'd0}, _T_2776}; // @[PALU.scala 428:38]
  wire [2:0] _T_2804 = _T_2803 + _GEN_655; // @[PALU.scala 428:38]
  wire [2:0] _GEN_656 = {{2'd0}, _T_2778}; // @[PALU.scala 428:38]
  wire [3:0] _T_2805 = _T_2804 + _GEN_656; // @[PALU.scala 428:38]
  wire [3:0] _GEN_657 = {{3'd0}, _T_2780}; // @[PALU.scala 428:38]
  wire [4:0] _T_2806 = _T_2805 + _GEN_657; // @[PALU.scala 428:38]
  wire [4:0] _GEN_658 = {{4'd0}, _T_2782}; // @[PALU.scala 428:38]
  wire [5:0] _T_2807 = _T_2806 + _GEN_658; // @[PALU.scala 428:38]
  wire [5:0] _GEN_659 = {{5'd0}, _T_2784}; // @[PALU.scala 428:38]
  wire [6:0] _T_2808 = _T_2807 + _GEN_659; // @[PALU.scala 428:38]
  wire [6:0] _GEN_660 = {{6'd0}, _T_2786}; // @[PALU.scala 428:38]
  wire [7:0] _T_2809 = _T_2808 + _GEN_660; // @[PALU.scala 428:38]
  wire [7:0] _GEN_661 = {{7'd0}, _T_2788}; // @[PALU.scala 428:38]
  wire [8:0] _T_2810 = _T_2809 + _GEN_661; // @[PALU.scala 428:38]
  wire [8:0] _GEN_662 = {{8'd0}, _T_2790}; // @[PALU.scala 428:38]
  wire [9:0] _T_2811 = _T_2810 + _GEN_662; // @[PALU.scala 428:38]
  wire [9:0] _GEN_663 = {{9'd0}, _T_2792}; // @[PALU.scala 428:38]
  wire [10:0] _T_2812 = _T_2811 + _GEN_663; // @[PALU.scala 428:38]
  wire [10:0] _GEN_664 = {{10'd0}, _T_2794}; // @[PALU.scala 428:38]
  wire [11:0] _T_2813 = _T_2812 + _GEN_664; // @[PALU.scala 428:38]
  wire [11:0] _GEN_665 = {{11'd0}, _T_2796}; // @[PALU.scala 428:38]
  wire [12:0] _T_2814 = _T_2813 + _GEN_665; // @[PALU.scala 428:38]
  wire [12:0] _GEN_666 = {{12'd0}, _T_2798}; // @[PALU.scala 428:38]
  wire [13:0] _T_2815 = _T_2814 + _GEN_666; // @[PALU.scala 428:38]
  wire [13:0] _GEN_667 = {{13'd0}, _T_2800}; // @[PALU.scala 428:38]
  wire [14:0] _T_2816 = _T_2815 + _GEN_667; // @[PALU.scala 428:38]
  wire [14:0] _GEN_668 = {{14'd0}, _T_2802}; // @[PALU.scala 428:38]
  wire [15:0] _T_2817 = _T_2816 + _GEN_668; // @[PALU.scala 428:38]
  wire [15:0] _T_2819 = _T_2817 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_2820 = io_in_bits_DecodeIn_data_src2[0] ? _T_2817 : _T_2819; // @[PALU.scala 429:26]
  wire  _T_2823 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[31]; // @[PALU.scala 423:29]
  wire  _T_2825 = io_in_bits_DecodeIn_data_src1[16] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2827 = io_in_bits_DecodeIn_data_src1[17] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2829 = io_in_bits_DecodeIn_data_src1[18] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2831 = io_in_bits_DecodeIn_data_src1[19] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2833 = io_in_bits_DecodeIn_data_src1[20] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2835 = io_in_bits_DecodeIn_data_src1[21] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2837 = io_in_bits_DecodeIn_data_src1[22] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2839 = io_in_bits_DecodeIn_data_src1[23] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2841 = io_in_bits_DecodeIn_data_src1[24] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2843 = io_in_bits_DecodeIn_data_src1[25] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2845 = io_in_bits_DecodeIn_data_src1[26] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2847 = io_in_bits_DecodeIn_data_src1[27] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2849 = io_in_bits_DecodeIn_data_src1[28] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2851 = io_in_bits_DecodeIn_data_src1[29] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2853 = io_in_bits_DecodeIn_data_src1[30] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2855 = io_in_bits_DecodeIn_data_src1[31] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2857 = _T_2853 & _T_2855; // @[PALU.scala 427:113]
  wire  _T_2859 = _T_2851 & (_T_2853 & _T_2855); // @[PALU.scala 427:113]
  wire  _T_2861 = _T_2849 & (_T_2851 & (_T_2853 & _T_2855)); // @[PALU.scala 427:113]
  wire  _T_2863 = _T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))); // @[PALU.scala 427:113]
  wire  _T_2865 = _T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))); // @[PALU.scala 427:113]
  wire  _T_2867 = _T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))))); // @[PALU.scala 427:113]
  wire  _T_2869 = _T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))))); // @[PALU.scala 427:113]
  wire  _T_2871 = _T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))))))); // @[PALU.scala 427:113]
  wire  _T_2873 = _T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 &
    _T_2855)))))))); // @[PALU.scala 427:113]
  wire  _T_2875 = _T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (
    _T_2853 & _T_2855))))))))); // @[PALU.scala 427:113]
  wire  _T_2877 = _T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (
    _T_2851 & (_T_2853 & _T_2855)))))))))); // @[PALU.scala 427:113]
  wire  _T_2879 = _T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (
    _T_2849 & (_T_2851 & (_T_2853 & _T_2855))))))))))); // @[PALU.scala 427:113]
  wire  _T_2881 = _T_2829 & (_T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (
    _T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))))))))))); // @[PALU.scala 427:113]
  wire  _T_2883 = _T_2827 & (_T_2829 & (_T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (
    _T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))))))))))))); // @[PALU.scala 427:113]
  wire  _T_2885 = _T_2825 & (_T_2827 & (_T_2829 & (_T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (
    _T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_2886 = _T_2855 + _T_2857; // @[PALU.scala 428:38]
  wire [1:0] _GEN_669 = {{1'd0}, _T_2859}; // @[PALU.scala 428:38]
  wire [2:0] _T_2887 = _T_2886 + _GEN_669; // @[PALU.scala 428:38]
  wire [2:0] _GEN_670 = {{2'd0}, _T_2861}; // @[PALU.scala 428:38]
  wire [3:0] _T_2888 = _T_2887 + _GEN_670; // @[PALU.scala 428:38]
  wire [3:0] _GEN_671 = {{3'd0}, _T_2863}; // @[PALU.scala 428:38]
  wire [4:0] _T_2889 = _T_2888 + _GEN_671; // @[PALU.scala 428:38]
  wire [4:0] _GEN_672 = {{4'd0}, _T_2865}; // @[PALU.scala 428:38]
  wire [5:0] _T_2890 = _T_2889 + _GEN_672; // @[PALU.scala 428:38]
  wire [5:0] _GEN_673 = {{5'd0}, _T_2867}; // @[PALU.scala 428:38]
  wire [6:0] _T_2891 = _T_2890 + _GEN_673; // @[PALU.scala 428:38]
  wire [6:0] _GEN_674 = {{6'd0}, _T_2869}; // @[PALU.scala 428:38]
  wire [7:0] _T_2892 = _T_2891 + _GEN_674; // @[PALU.scala 428:38]
  wire [7:0] _GEN_675 = {{7'd0}, _T_2871}; // @[PALU.scala 428:38]
  wire [8:0] _T_2893 = _T_2892 + _GEN_675; // @[PALU.scala 428:38]
  wire [8:0] _GEN_676 = {{8'd0}, _T_2873}; // @[PALU.scala 428:38]
  wire [9:0] _T_2894 = _T_2893 + _GEN_676; // @[PALU.scala 428:38]
  wire [9:0] _GEN_677 = {{9'd0}, _T_2875}; // @[PALU.scala 428:38]
  wire [10:0] _T_2895 = _T_2894 + _GEN_677; // @[PALU.scala 428:38]
  wire [10:0] _GEN_678 = {{10'd0}, _T_2877}; // @[PALU.scala 428:38]
  wire [11:0] _T_2896 = _T_2895 + _GEN_678; // @[PALU.scala 428:38]
  wire [11:0] _GEN_679 = {{11'd0}, _T_2879}; // @[PALU.scala 428:38]
  wire [12:0] _T_2897 = _T_2896 + _GEN_679; // @[PALU.scala 428:38]
  wire [12:0] _GEN_680 = {{12'd0}, _T_2881}; // @[PALU.scala 428:38]
  wire [13:0] _T_2898 = _T_2897 + _GEN_680; // @[PALU.scala 428:38]
  wire [13:0] _GEN_681 = {{13'd0}, _T_2883}; // @[PALU.scala 428:38]
  wire [14:0] _T_2899 = _T_2898 + _GEN_681; // @[PALU.scala 428:38]
  wire [14:0] _GEN_682 = {{14'd0}, _T_2885}; // @[PALU.scala 428:38]
  wire [15:0] _T_2900 = _T_2899 + _GEN_682; // @[PALU.scala 428:38]
  wire [15:0] _T_2902 = _T_2900 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_2903 = io_in_bits_DecodeIn_data_src2[0] ? _T_2900 : _T_2902; // @[PALU.scala 429:26]
  wire  _T_2906 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[47]; // @[PALU.scala 423:29]
  wire  _T_2908 = io_in_bits_DecodeIn_data_src1[32] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2910 = io_in_bits_DecodeIn_data_src1[33] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2912 = io_in_bits_DecodeIn_data_src1[34] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2914 = io_in_bits_DecodeIn_data_src1[35] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2916 = io_in_bits_DecodeIn_data_src1[36] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2918 = io_in_bits_DecodeIn_data_src1[37] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2920 = io_in_bits_DecodeIn_data_src1[38] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2922 = io_in_bits_DecodeIn_data_src1[39] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2924 = io_in_bits_DecodeIn_data_src1[40] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2926 = io_in_bits_DecodeIn_data_src1[41] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2928 = io_in_bits_DecodeIn_data_src1[42] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2930 = io_in_bits_DecodeIn_data_src1[43] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2932 = io_in_bits_DecodeIn_data_src1[44] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2934 = io_in_bits_DecodeIn_data_src1[45] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2936 = io_in_bits_DecodeIn_data_src1[46] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2938 = io_in_bits_DecodeIn_data_src1[47] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2940 = _T_2936 & _T_2938; // @[PALU.scala 427:113]
  wire  _T_2942 = _T_2934 & (_T_2936 & _T_2938); // @[PALU.scala 427:113]
  wire  _T_2944 = _T_2932 & (_T_2934 & (_T_2936 & _T_2938)); // @[PALU.scala 427:113]
  wire  _T_2946 = _T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))); // @[PALU.scala 427:113]
  wire  _T_2948 = _T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))); // @[PALU.scala 427:113]
  wire  _T_2950 = _T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))))); // @[PALU.scala 427:113]
  wire  _T_2952 = _T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))))); // @[PALU.scala 427:113]
  wire  _T_2954 = _T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))))))); // @[PALU.scala 427:113]
  wire  _T_2956 = _T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 &
    _T_2938)))))))); // @[PALU.scala 427:113]
  wire  _T_2958 = _T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (
    _T_2936 & _T_2938))))))))); // @[PALU.scala 427:113]
  wire  _T_2960 = _T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (
    _T_2934 & (_T_2936 & _T_2938)))))))))); // @[PALU.scala 427:113]
  wire  _T_2962 = _T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (
    _T_2932 & (_T_2934 & (_T_2936 & _T_2938))))))))))); // @[PALU.scala 427:113]
  wire  _T_2964 = _T_2912 & (_T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (
    _T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))))))))))); // @[PALU.scala 427:113]
  wire  _T_2966 = _T_2910 & (_T_2912 & (_T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (
    _T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))))))))))))); // @[PALU.scala 427:113]
  wire  _T_2968 = _T_2908 & (_T_2910 & (_T_2912 & (_T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (
    _T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_2969 = _T_2938 + _T_2940; // @[PALU.scala 428:38]
  wire [1:0] _GEN_683 = {{1'd0}, _T_2942}; // @[PALU.scala 428:38]
  wire [2:0] _T_2970 = _T_2969 + _GEN_683; // @[PALU.scala 428:38]
  wire [2:0] _GEN_684 = {{2'd0}, _T_2944}; // @[PALU.scala 428:38]
  wire [3:0] _T_2971 = _T_2970 + _GEN_684; // @[PALU.scala 428:38]
  wire [3:0] _GEN_685 = {{3'd0}, _T_2946}; // @[PALU.scala 428:38]
  wire [4:0] _T_2972 = _T_2971 + _GEN_685; // @[PALU.scala 428:38]
  wire [4:0] _GEN_686 = {{4'd0}, _T_2948}; // @[PALU.scala 428:38]
  wire [5:0] _T_2973 = _T_2972 + _GEN_686; // @[PALU.scala 428:38]
  wire [5:0] _GEN_687 = {{5'd0}, _T_2950}; // @[PALU.scala 428:38]
  wire [6:0] _T_2974 = _T_2973 + _GEN_687; // @[PALU.scala 428:38]
  wire [6:0] _GEN_688 = {{6'd0}, _T_2952}; // @[PALU.scala 428:38]
  wire [7:0] _T_2975 = _T_2974 + _GEN_688; // @[PALU.scala 428:38]
  wire [7:0] _GEN_689 = {{7'd0}, _T_2954}; // @[PALU.scala 428:38]
  wire [8:0] _T_2976 = _T_2975 + _GEN_689; // @[PALU.scala 428:38]
  wire [8:0] _GEN_690 = {{8'd0}, _T_2956}; // @[PALU.scala 428:38]
  wire [9:0] _T_2977 = _T_2976 + _GEN_690; // @[PALU.scala 428:38]
  wire [9:0] _GEN_691 = {{9'd0}, _T_2958}; // @[PALU.scala 428:38]
  wire [10:0] _T_2978 = _T_2977 + _GEN_691; // @[PALU.scala 428:38]
  wire [10:0] _GEN_692 = {{10'd0}, _T_2960}; // @[PALU.scala 428:38]
  wire [11:0] _T_2979 = _T_2978 + _GEN_692; // @[PALU.scala 428:38]
  wire [11:0] _GEN_693 = {{11'd0}, _T_2962}; // @[PALU.scala 428:38]
  wire [12:0] _T_2980 = _T_2979 + _GEN_693; // @[PALU.scala 428:38]
  wire [12:0] _GEN_694 = {{12'd0}, _T_2964}; // @[PALU.scala 428:38]
  wire [13:0] _T_2981 = _T_2980 + _GEN_694; // @[PALU.scala 428:38]
  wire [13:0] _GEN_695 = {{13'd0}, _T_2966}; // @[PALU.scala 428:38]
  wire [14:0] _T_2982 = _T_2981 + _GEN_695; // @[PALU.scala 428:38]
  wire [14:0] _GEN_696 = {{14'd0}, _T_2968}; // @[PALU.scala 428:38]
  wire [15:0] _T_2983 = _T_2982 + _GEN_696; // @[PALU.scala 428:38]
  wire [15:0] _T_2985 = _T_2983 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_2986 = io_in_bits_DecodeIn_data_src2[0] ? _T_2983 : _T_2985; // @[PALU.scala 429:26]
  wire  _T_2989 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[63]; // @[PALU.scala 423:29]
  wire  _T_2991 = io_in_bits_DecodeIn_data_src1[48] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2993 = io_in_bits_DecodeIn_data_src1[49] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2995 = io_in_bits_DecodeIn_data_src1[50] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2997 = io_in_bits_DecodeIn_data_src1[51] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2999 = io_in_bits_DecodeIn_data_src1[52] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3001 = io_in_bits_DecodeIn_data_src1[53] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3003 = io_in_bits_DecodeIn_data_src1[54] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3005 = io_in_bits_DecodeIn_data_src1[55] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3007 = io_in_bits_DecodeIn_data_src1[56] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3009 = io_in_bits_DecodeIn_data_src1[57] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3011 = io_in_bits_DecodeIn_data_src1[58] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3013 = io_in_bits_DecodeIn_data_src1[59] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3015 = io_in_bits_DecodeIn_data_src1[60] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3017 = io_in_bits_DecodeIn_data_src1[61] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3019 = io_in_bits_DecodeIn_data_src1[62] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3021 = io_in_bits_DecodeIn_data_src1[63] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3023 = _T_3019 & _T_3021; // @[PALU.scala 427:113]
  wire  _T_3025 = _T_3017 & (_T_3019 & _T_3021); // @[PALU.scala 427:113]
  wire  _T_3027 = _T_3015 & (_T_3017 & (_T_3019 & _T_3021)); // @[PALU.scala 427:113]
  wire  _T_3029 = _T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))); // @[PALU.scala 427:113]
  wire  _T_3031 = _T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))); // @[PALU.scala 427:113]
  wire  _T_3033 = _T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))))); // @[PALU.scala 427:113]
  wire  _T_3035 = _T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))))); // @[PALU.scala 427:113]
  wire  _T_3037 = _T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))))))); // @[PALU.scala 427:113]
  wire  _T_3039 = _T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 &
    _T_3021)))))))); // @[PALU.scala 427:113]
  wire  _T_3041 = _T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (
    _T_3019 & _T_3021))))))))); // @[PALU.scala 427:113]
  wire  _T_3043 = _T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (
    _T_3017 & (_T_3019 & _T_3021)))))))))); // @[PALU.scala 427:113]
  wire  _T_3045 = _T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (
    _T_3015 & (_T_3017 & (_T_3019 & _T_3021))))))))))); // @[PALU.scala 427:113]
  wire  _T_3047 = _T_2995 & (_T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (
    _T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))))))))))); // @[PALU.scala 427:113]
  wire  _T_3049 = _T_2993 & (_T_2995 & (_T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (
    _T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3051 = _T_2991 & (_T_2993 & (_T_2995 & (_T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (
    _T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3052 = _T_3021 + _T_3023; // @[PALU.scala 428:38]
  wire [1:0] _GEN_697 = {{1'd0}, _T_3025}; // @[PALU.scala 428:38]
  wire [2:0] _T_3053 = _T_3052 + _GEN_697; // @[PALU.scala 428:38]
  wire [2:0] _GEN_698 = {{2'd0}, _T_3027}; // @[PALU.scala 428:38]
  wire [3:0] _T_3054 = _T_3053 + _GEN_698; // @[PALU.scala 428:38]
  wire [3:0] _GEN_699 = {{3'd0}, _T_3029}; // @[PALU.scala 428:38]
  wire [4:0] _T_3055 = _T_3054 + _GEN_699; // @[PALU.scala 428:38]
  wire [4:0] _GEN_700 = {{4'd0}, _T_3031}; // @[PALU.scala 428:38]
  wire [5:0] _T_3056 = _T_3055 + _GEN_700; // @[PALU.scala 428:38]
  wire [5:0] _GEN_701 = {{5'd0}, _T_3033}; // @[PALU.scala 428:38]
  wire [6:0] _T_3057 = _T_3056 + _GEN_701; // @[PALU.scala 428:38]
  wire [6:0] _GEN_702 = {{6'd0}, _T_3035}; // @[PALU.scala 428:38]
  wire [7:0] _T_3058 = _T_3057 + _GEN_702; // @[PALU.scala 428:38]
  wire [7:0] _GEN_703 = {{7'd0}, _T_3037}; // @[PALU.scala 428:38]
  wire [8:0] _T_3059 = _T_3058 + _GEN_703; // @[PALU.scala 428:38]
  wire [8:0] _GEN_704 = {{8'd0}, _T_3039}; // @[PALU.scala 428:38]
  wire [9:0] _T_3060 = _T_3059 + _GEN_704; // @[PALU.scala 428:38]
  wire [9:0] _GEN_705 = {{9'd0}, _T_3041}; // @[PALU.scala 428:38]
  wire [10:0] _T_3061 = _T_3060 + _GEN_705; // @[PALU.scala 428:38]
  wire [10:0] _GEN_706 = {{10'd0}, _T_3043}; // @[PALU.scala 428:38]
  wire [11:0] _T_3062 = _T_3061 + _GEN_706; // @[PALU.scala 428:38]
  wire [11:0] _GEN_707 = {{11'd0}, _T_3045}; // @[PALU.scala 428:38]
  wire [12:0] _T_3063 = _T_3062 + _GEN_707; // @[PALU.scala 428:38]
  wire [12:0] _GEN_708 = {{12'd0}, _T_3047}; // @[PALU.scala 428:38]
  wire [13:0] _T_3064 = _T_3063 + _GEN_708; // @[PALU.scala 428:38]
  wire [13:0] _GEN_709 = {{13'd0}, _T_3049}; // @[PALU.scala 428:38]
  wire [14:0] _T_3065 = _T_3064 + _GEN_709; // @[PALU.scala 428:38]
  wire [14:0] _GEN_710 = {{14'd0}, _T_3051}; // @[PALU.scala 428:38]
  wire [15:0] _T_3066 = _T_3065 + _GEN_710; // @[PALU.scala 428:38]
  wire [15:0] _T_3068 = _T_3066 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_3069 = io_in_bits_DecodeIn_data_src2[0] ? _T_3066 : _T_3068; // @[PALU.scala 429:26]
  wire [63:0] _T_3072 = {_T_3069,_T_2986,_T_2903,_T_2820}; // @[Cat.scala 30:58]
  wire  _T_3077 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[7]; // @[PALU.scala 423:29]
  wire  _T_3079 = io_in_bits_DecodeIn_data_src1[0] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3081 = io_in_bits_DecodeIn_data_src1[1] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3083 = io_in_bits_DecodeIn_data_src1[2] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3085 = io_in_bits_DecodeIn_data_src1[3] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3087 = io_in_bits_DecodeIn_data_src1[4] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3089 = io_in_bits_DecodeIn_data_src1[5] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3091 = io_in_bits_DecodeIn_data_src1[6] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3093 = io_in_bits_DecodeIn_data_src1[7] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3095 = _T_3091 & _T_3093; // @[PALU.scala 427:113]
  wire  _T_3097 = _T_3089 & (_T_3091 & _T_3093); // @[PALU.scala 427:113]
  wire  _T_3099 = _T_3087 & (_T_3089 & (_T_3091 & _T_3093)); // @[PALU.scala 427:113]
  wire  _T_3101 = _T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093))); // @[PALU.scala 427:113]
  wire  _T_3103 = _T_3083 & (_T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093)))); // @[PALU.scala 427:113]
  wire  _T_3105 = _T_3081 & (_T_3083 & (_T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093))))); // @[PALU.scala 427:113]
  wire  _T_3107 = _T_3079 & (_T_3081 & (_T_3083 & (_T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3108 = _T_3093 + _T_3095; // @[PALU.scala 428:38]
  wire [1:0] _GEN_711 = {{1'd0}, _T_3097}; // @[PALU.scala 428:38]
  wire [2:0] _T_3109 = _T_3108 + _GEN_711; // @[PALU.scala 428:38]
  wire [2:0] _GEN_712 = {{2'd0}, _T_3099}; // @[PALU.scala 428:38]
  wire [3:0] _T_3110 = _T_3109 + _GEN_712; // @[PALU.scala 428:38]
  wire [3:0] _GEN_713 = {{3'd0}, _T_3101}; // @[PALU.scala 428:38]
  wire [4:0] _T_3111 = _T_3110 + _GEN_713; // @[PALU.scala 428:38]
  wire [4:0] _GEN_714 = {{4'd0}, _T_3103}; // @[PALU.scala 428:38]
  wire [5:0] _T_3112 = _T_3111 + _GEN_714; // @[PALU.scala 428:38]
  wire [5:0] _GEN_715 = {{5'd0}, _T_3105}; // @[PALU.scala 428:38]
  wire [6:0] _T_3113 = _T_3112 + _GEN_715; // @[PALU.scala 428:38]
  wire [6:0] _GEN_716 = {{6'd0}, _T_3107}; // @[PALU.scala 428:38]
  wire [7:0] _T_3114 = _T_3113 + _GEN_716; // @[PALU.scala 428:38]
  wire [7:0] _T_3116 = _T_3114 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3117 = io_in_bits_DecodeIn_data_src2[0] ? _T_3114 : _T_3116; // @[PALU.scala 429:26]
  wire  _T_3120 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[15]; // @[PALU.scala 423:29]
  wire  _T_3122 = io_in_bits_DecodeIn_data_src1[8] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3124 = io_in_bits_DecodeIn_data_src1[9] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3126 = io_in_bits_DecodeIn_data_src1[10] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3128 = io_in_bits_DecodeIn_data_src1[11] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3130 = io_in_bits_DecodeIn_data_src1[12] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3132 = io_in_bits_DecodeIn_data_src1[13] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3134 = io_in_bits_DecodeIn_data_src1[14] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3136 = io_in_bits_DecodeIn_data_src1[15] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3138 = _T_3134 & _T_3136; // @[PALU.scala 427:113]
  wire  _T_3140 = _T_3132 & (_T_3134 & _T_3136); // @[PALU.scala 427:113]
  wire  _T_3142 = _T_3130 & (_T_3132 & (_T_3134 & _T_3136)); // @[PALU.scala 427:113]
  wire  _T_3144 = _T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136))); // @[PALU.scala 427:113]
  wire  _T_3146 = _T_3126 & (_T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136)))); // @[PALU.scala 427:113]
  wire  _T_3148 = _T_3124 & (_T_3126 & (_T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136))))); // @[PALU.scala 427:113]
  wire  _T_3150 = _T_3122 & (_T_3124 & (_T_3126 & (_T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3151 = _T_3136 + _T_3138; // @[PALU.scala 428:38]
  wire [1:0] _GEN_717 = {{1'd0}, _T_3140}; // @[PALU.scala 428:38]
  wire [2:0] _T_3152 = _T_3151 + _GEN_717; // @[PALU.scala 428:38]
  wire [2:0] _GEN_718 = {{2'd0}, _T_3142}; // @[PALU.scala 428:38]
  wire [3:0] _T_3153 = _T_3152 + _GEN_718; // @[PALU.scala 428:38]
  wire [3:0] _GEN_719 = {{3'd0}, _T_3144}; // @[PALU.scala 428:38]
  wire [4:0] _T_3154 = _T_3153 + _GEN_719; // @[PALU.scala 428:38]
  wire [4:0] _GEN_720 = {{4'd0}, _T_3146}; // @[PALU.scala 428:38]
  wire [5:0] _T_3155 = _T_3154 + _GEN_720; // @[PALU.scala 428:38]
  wire [5:0] _GEN_721 = {{5'd0}, _T_3148}; // @[PALU.scala 428:38]
  wire [6:0] _T_3156 = _T_3155 + _GEN_721; // @[PALU.scala 428:38]
  wire [6:0] _GEN_722 = {{6'd0}, _T_3150}; // @[PALU.scala 428:38]
  wire [7:0] _T_3157 = _T_3156 + _GEN_722; // @[PALU.scala 428:38]
  wire [7:0] _T_3159 = _T_3157 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3160 = io_in_bits_DecodeIn_data_src2[0] ? _T_3157 : _T_3159; // @[PALU.scala 429:26]
  wire  _T_3163 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[23]; // @[PALU.scala 423:29]
  wire  _T_3165 = io_in_bits_DecodeIn_data_src1[16] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3167 = io_in_bits_DecodeIn_data_src1[17] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3169 = io_in_bits_DecodeIn_data_src1[18] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3171 = io_in_bits_DecodeIn_data_src1[19] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3173 = io_in_bits_DecodeIn_data_src1[20] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3175 = io_in_bits_DecodeIn_data_src1[21] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3177 = io_in_bits_DecodeIn_data_src1[22] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3179 = io_in_bits_DecodeIn_data_src1[23] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3181 = _T_3177 & _T_3179; // @[PALU.scala 427:113]
  wire  _T_3183 = _T_3175 & (_T_3177 & _T_3179); // @[PALU.scala 427:113]
  wire  _T_3185 = _T_3173 & (_T_3175 & (_T_3177 & _T_3179)); // @[PALU.scala 427:113]
  wire  _T_3187 = _T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179))); // @[PALU.scala 427:113]
  wire  _T_3189 = _T_3169 & (_T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179)))); // @[PALU.scala 427:113]
  wire  _T_3191 = _T_3167 & (_T_3169 & (_T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179))))); // @[PALU.scala 427:113]
  wire  _T_3193 = _T_3165 & (_T_3167 & (_T_3169 & (_T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3194 = _T_3179 + _T_3181; // @[PALU.scala 428:38]
  wire [1:0] _GEN_723 = {{1'd0}, _T_3183}; // @[PALU.scala 428:38]
  wire [2:0] _T_3195 = _T_3194 + _GEN_723; // @[PALU.scala 428:38]
  wire [2:0] _GEN_724 = {{2'd0}, _T_3185}; // @[PALU.scala 428:38]
  wire [3:0] _T_3196 = _T_3195 + _GEN_724; // @[PALU.scala 428:38]
  wire [3:0] _GEN_725 = {{3'd0}, _T_3187}; // @[PALU.scala 428:38]
  wire [4:0] _T_3197 = _T_3196 + _GEN_725; // @[PALU.scala 428:38]
  wire [4:0] _GEN_726 = {{4'd0}, _T_3189}; // @[PALU.scala 428:38]
  wire [5:0] _T_3198 = _T_3197 + _GEN_726; // @[PALU.scala 428:38]
  wire [5:0] _GEN_727 = {{5'd0}, _T_3191}; // @[PALU.scala 428:38]
  wire [6:0] _T_3199 = _T_3198 + _GEN_727; // @[PALU.scala 428:38]
  wire [6:0] _GEN_728 = {{6'd0}, _T_3193}; // @[PALU.scala 428:38]
  wire [7:0] _T_3200 = _T_3199 + _GEN_728; // @[PALU.scala 428:38]
  wire [7:0] _T_3202 = _T_3200 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3203 = io_in_bits_DecodeIn_data_src2[0] ? _T_3200 : _T_3202; // @[PALU.scala 429:26]
  wire  _T_3206 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[31]; // @[PALU.scala 423:29]
  wire  _T_3208 = io_in_bits_DecodeIn_data_src1[24] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3210 = io_in_bits_DecodeIn_data_src1[25] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3212 = io_in_bits_DecodeIn_data_src1[26] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3214 = io_in_bits_DecodeIn_data_src1[27] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3216 = io_in_bits_DecodeIn_data_src1[28] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3218 = io_in_bits_DecodeIn_data_src1[29] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3220 = io_in_bits_DecodeIn_data_src1[30] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3222 = io_in_bits_DecodeIn_data_src1[31] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3224 = _T_3220 & _T_3222; // @[PALU.scala 427:113]
  wire  _T_3226 = _T_3218 & (_T_3220 & _T_3222); // @[PALU.scala 427:113]
  wire  _T_3228 = _T_3216 & (_T_3218 & (_T_3220 & _T_3222)); // @[PALU.scala 427:113]
  wire  _T_3230 = _T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222))); // @[PALU.scala 427:113]
  wire  _T_3232 = _T_3212 & (_T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222)))); // @[PALU.scala 427:113]
  wire  _T_3234 = _T_3210 & (_T_3212 & (_T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222))))); // @[PALU.scala 427:113]
  wire  _T_3236 = _T_3208 & (_T_3210 & (_T_3212 & (_T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3237 = _T_3222 + _T_3224; // @[PALU.scala 428:38]
  wire [1:0] _GEN_729 = {{1'd0}, _T_3226}; // @[PALU.scala 428:38]
  wire [2:0] _T_3238 = _T_3237 + _GEN_729; // @[PALU.scala 428:38]
  wire [2:0] _GEN_730 = {{2'd0}, _T_3228}; // @[PALU.scala 428:38]
  wire [3:0] _T_3239 = _T_3238 + _GEN_730; // @[PALU.scala 428:38]
  wire [3:0] _GEN_731 = {{3'd0}, _T_3230}; // @[PALU.scala 428:38]
  wire [4:0] _T_3240 = _T_3239 + _GEN_731; // @[PALU.scala 428:38]
  wire [4:0] _GEN_732 = {{4'd0}, _T_3232}; // @[PALU.scala 428:38]
  wire [5:0] _T_3241 = _T_3240 + _GEN_732; // @[PALU.scala 428:38]
  wire [5:0] _GEN_733 = {{5'd0}, _T_3234}; // @[PALU.scala 428:38]
  wire [6:0] _T_3242 = _T_3241 + _GEN_733; // @[PALU.scala 428:38]
  wire [6:0] _GEN_734 = {{6'd0}, _T_3236}; // @[PALU.scala 428:38]
  wire [7:0] _T_3243 = _T_3242 + _GEN_734; // @[PALU.scala 428:38]
  wire [7:0] _T_3245 = _T_3243 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3246 = io_in_bits_DecodeIn_data_src2[0] ? _T_3243 : _T_3245; // @[PALU.scala 429:26]
  wire  _T_3249 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[39]; // @[PALU.scala 423:29]
  wire  _T_3251 = io_in_bits_DecodeIn_data_src1[32] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3253 = io_in_bits_DecodeIn_data_src1[33] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3255 = io_in_bits_DecodeIn_data_src1[34] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3257 = io_in_bits_DecodeIn_data_src1[35] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3259 = io_in_bits_DecodeIn_data_src1[36] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3261 = io_in_bits_DecodeIn_data_src1[37] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3263 = io_in_bits_DecodeIn_data_src1[38] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3265 = io_in_bits_DecodeIn_data_src1[39] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3267 = _T_3263 & _T_3265; // @[PALU.scala 427:113]
  wire  _T_3269 = _T_3261 & (_T_3263 & _T_3265); // @[PALU.scala 427:113]
  wire  _T_3271 = _T_3259 & (_T_3261 & (_T_3263 & _T_3265)); // @[PALU.scala 427:113]
  wire  _T_3273 = _T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265))); // @[PALU.scala 427:113]
  wire  _T_3275 = _T_3255 & (_T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265)))); // @[PALU.scala 427:113]
  wire  _T_3277 = _T_3253 & (_T_3255 & (_T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265))))); // @[PALU.scala 427:113]
  wire  _T_3279 = _T_3251 & (_T_3253 & (_T_3255 & (_T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3280 = _T_3265 + _T_3267; // @[PALU.scala 428:38]
  wire [1:0] _GEN_735 = {{1'd0}, _T_3269}; // @[PALU.scala 428:38]
  wire [2:0] _T_3281 = _T_3280 + _GEN_735; // @[PALU.scala 428:38]
  wire [2:0] _GEN_736 = {{2'd0}, _T_3271}; // @[PALU.scala 428:38]
  wire [3:0] _T_3282 = _T_3281 + _GEN_736; // @[PALU.scala 428:38]
  wire [3:0] _GEN_737 = {{3'd0}, _T_3273}; // @[PALU.scala 428:38]
  wire [4:0] _T_3283 = _T_3282 + _GEN_737; // @[PALU.scala 428:38]
  wire [4:0] _GEN_738 = {{4'd0}, _T_3275}; // @[PALU.scala 428:38]
  wire [5:0] _T_3284 = _T_3283 + _GEN_738; // @[PALU.scala 428:38]
  wire [5:0] _GEN_739 = {{5'd0}, _T_3277}; // @[PALU.scala 428:38]
  wire [6:0] _T_3285 = _T_3284 + _GEN_739; // @[PALU.scala 428:38]
  wire [6:0] _GEN_740 = {{6'd0}, _T_3279}; // @[PALU.scala 428:38]
  wire [7:0] _T_3286 = _T_3285 + _GEN_740; // @[PALU.scala 428:38]
  wire [7:0] _T_3288 = _T_3286 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3289 = io_in_bits_DecodeIn_data_src2[0] ? _T_3286 : _T_3288; // @[PALU.scala 429:26]
  wire  _T_3292 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[47]; // @[PALU.scala 423:29]
  wire  _T_3294 = io_in_bits_DecodeIn_data_src1[40] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3296 = io_in_bits_DecodeIn_data_src1[41] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3298 = io_in_bits_DecodeIn_data_src1[42] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3300 = io_in_bits_DecodeIn_data_src1[43] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3302 = io_in_bits_DecodeIn_data_src1[44] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3304 = io_in_bits_DecodeIn_data_src1[45] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3306 = io_in_bits_DecodeIn_data_src1[46] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3308 = io_in_bits_DecodeIn_data_src1[47] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3310 = _T_3306 & _T_3308; // @[PALU.scala 427:113]
  wire  _T_3312 = _T_3304 & (_T_3306 & _T_3308); // @[PALU.scala 427:113]
  wire  _T_3314 = _T_3302 & (_T_3304 & (_T_3306 & _T_3308)); // @[PALU.scala 427:113]
  wire  _T_3316 = _T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308))); // @[PALU.scala 427:113]
  wire  _T_3318 = _T_3298 & (_T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308)))); // @[PALU.scala 427:113]
  wire  _T_3320 = _T_3296 & (_T_3298 & (_T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308))))); // @[PALU.scala 427:113]
  wire  _T_3322 = _T_3294 & (_T_3296 & (_T_3298 & (_T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3323 = _T_3308 + _T_3310; // @[PALU.scala 428:38]
  wire [1:0] _GEN_741 = {{1'd0}, _T_3312}; // @[PALU.scala 428:38]
  wire [2:0] _T_3324 = _T_3323 + _GEN_741; // @[PALU.scala 428:38]
  wire [2:0] _GEN_742 = {{2'd0}, _T_3314}; // @[PALU.scala 428:38]
  wire [3:0] _T_3325 = _T_3324 + _GEN_742; // @[PALU.scala 428:38]
  wire [3:0] _GEN_743 = {{3'd0}, _T_3316}; // @[PALU.scala 428:38]
  wire [4:0] _T_3326 = _T_3325 + _GEN_743; // @[PALU.scala 428:38]
  wire [4:0] _GEN_744 = {{4'd0}, _T_3318}; // @[PALU.scala 428:38]
  wire [5:0] _T_3327 = _T_3326 + _GEN_744; // @[PALU.scala 428:38]
  wire [5:0] _GEN_745 = {{5'd0}, _T_3320}; // @[PALU.scala 428:38]
  wire [6:0] _T_3328 = _T_3327 + _GEN_745; // @[PALU.scala 428:38]
  wire [6:0] _GEN_746 = {{6'd0}, _T_3322}; // @[PALU.scala 428:38]
  wire [7:0] _T_3329 = _T_3328 + _GEN_746; // @[PALU.scala 428:38]
  wire [7:0] _T_3331 = _T_3329 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3332 = io_in_bits_DecodeIn_data_src2[0] ? _T_3329 : _T_3331; // @[PALU.scala 429:26]
  wire  _T_3335 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[55]; // @[PALU.scala 423:29]
  wire  _T_3337 = io_in_bits_DecodeIn_data_src1[48] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3339 = io_in_bits_DecodeIn_data_src1[49] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3341 = io_in_bits_DecodeIn_data_src1[50] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3343 = io_in_bits_DecodeIn_data_src1[51] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3345 = io_in_bits_DecodeIn_data_src1[52] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3347 = io_in_bits_DecodeIn_data_src1[53] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3349 = io_in_bits_DecodeIn_data_src1[54] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3351 = io_in_bits_DecodeIn_data_src1[55] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3353 = _T_3349 & _T_3351; // @[PALU.scala 427:113]
  wire  _T_3355 = _T_3347 & (_T_3349 & _T_3351); // @[PALU.scala 427:113]
  wire  _T_3357 = _T_3345 & (_T_3347 & (_T_3349 & _T_3351)); // @[PALU.scala 427:113]
  wire  _T_3359 = _T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351))); // @[PALU.scala 427:113]
  wire  _T_3361 = _T_3341 & (_T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351)))); // @[PALU.scala 427:113]
  wire  _T_3363 = _T_3339 & (_T_3341 & (_T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351))))); // @[PALU.scala 427:113]
  wire  _T_3365 = _T_3337 & (_T_3339 & (_T_3341 & (_T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3366 = _T_3351 + _T_3353; // @[PALU.scala 428:38]
  wire [1:0] _GEN_747 = {{1'd0}, _T_3355}; // @[PALU.scala 428:38]
  wire [2:0] _T_3367 = _T_3366 + _GEN_747; // @[PALU.scala 428:38]
  wire [2:0] _GEN_748 = {{2'd0}, _T_3357}; // @[PALU.scala 428:38]
  wire [3:0] _T_3368 = _T_3367 + _GEN_748; // @[PALU.scala 428:38]
  wire [3:0] _GEN_749 = {{3'd0}, _T_3359}; // @[PALU.scala 428:38]
  wire [4:0] _T_3369 = _T_3368 + _GEN_749; // @[PALU.scala 428:38]
  wire [4:0] _GEN_750 = {{4'd0}, _T_3361}; // @[PALU.scala 428:38]
  wire [5:0] _T_3370 = _T_3369 + _GEN_750; // @[PALU.scala 428:38]
  wire [5:0] _GEN_751 = {{5'd0}, _T_3363}; // @[PALU.scala 428:38]
  wire [6:0] _T_3371 = _T_3370 + _GEN_751; // @[PALU.scala 428:38]
  wire [6:0] _GEN_752 = {{6'd0}, _T_3365}; // @[PALU.scala 428:38]
  wire [7:0] _T_3372 = _T_3371 + _GEN_752; // @[PALU.scala 428:38]
  wire [7:0] _T_3374 = _T_3372 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3375 = io_in_bits_DecodeIn_data_src2[0] ? _T_3372 : _T_3374; // @[PALU.scala 429:26]
  wire  _T_3378 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[63]; // @[PALU.scala 423:29]
  wire  _T_3380 = io_in_bits_DecodeIn_data_src1[56] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3382 = io_in_bits_DecodeIn_data_src1[57] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3384 = io_in_bits_DecodeIn_data_src1[58] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3386 = io_in_bits_DecodeIn_data_src1[59] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3388 = io_in_bits_DecodeIn_data_src1[60] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3390 = io_in_bits_DecodeIn_data_src1[61] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3392 = io_in_bits_DecodeIn_data_src1[62] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3394 = io_in_bits_DecodeIn_data_src1[63] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3396 = _T_3392 & _T_3394; // @[PALU.scala 427:113]
  wire  _T_3398 = _T_3390 & (_T_3392 & _T_3394); // @[PALU.scala 427:113]
  wire  _T_3400 = _T_3388 & (_T_3390 & (_T_3392 & _T_3394)); // @[PALU.scala 427:113]
  wire  _T_3402 = _T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394))); // @[PALU.scala 427:113]
  wire  _T_3404 = _T_3384 & (_T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394)))); // @[PALU.scala 427:113]
  wire  _T_3406 = _T_3382 & (_T_3384 & (_T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394))))); // @[PALU.scala 427:113]
  wire  _T_3408 = _T_3380 & (_T_3382 & (_T_3384 & (_T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3409 = _T_3394 + _T_3396; // @[PALU.scala 428:38]
  wire [1:0] _GEN_753 = {{1'd0}, _T_3398}; // @[PALU.scala 428:38]
  wire [2:0] _T_3410 = _T_3409 + _GEN_753; // @[PALU.scala 428:38]
  wire [2:0] _GEN_754 = {{2'd0}, _T_3400}; // @[PALU.scala 428:38]
  wire [3:0] _T_3411 = _T_3410 + _GEN_754; // @[PALU.scala 428:38]
  wire [3:0] _GEN_755 = {{3'd0}, _T_3402}; // @[PALU.scala 428:38]
  wire [4:0] _T_3412 = _T_3411 + _GEN_755; // @[PALU.scala 428:38]
  wire [4:0] _GEN_756 = {{4'd0}, _T_3404}; // @[PALU.scala 428:38]
  wire [5:0] _T_3413 = _T_3412 + _GEN_756; // @[PALU.scala 428:38]
  wire [5:0] _GEN_757 = {{5'd0}, _T_3406}; // @[PALU.scala 428:38]
  wire [6:0] _T_3414 = _T_3413 + _GEN_757; // @[PALU.scala 428:38]
  wire [6:0] _GEN_758 = {{6'd0}, _T_3408}; // @[PALU.scala 428:38]
  wire [7:0] _T_3415 = _T_3414 + _GEN_758; // @[PALU.scala 428:38]
  wire [7:0] _T_3417 = _T_3415 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3418 = io_in_bits_DecodeIn_data_src2[0] ? _T_3415 : _T_3417; // @[PALU.scala 429:26]
  wire [63:0] _T_3425 = {_T_3418,_T_3375,_T_3332,_T_3289,_T_3246,_T_3203,_T_3160,_T_3117}; // @[Cat.scala 30:58]
  wire  _T_3430 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[31]; // @[PALU.scala 423:29]
  wire  _T_3432 = io_in_bits_DecodeIn_data_src1[0] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3434 = io_in_bits_DecodeIn_data_src1[1] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3436 = io_in_bits_DecodeIn_data_src1[2] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3438 = io_in_bits_DecodeIn_data_src1[3] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3440 = io_in_bits_DecodeIn_data_src1[4] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3442 = io_in_bits_DecodeIn_data_src1[5] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3444 = io_in_bits_DecodeIn_data_src1[6] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3446 = io_in_bits_DecodeIn_data_src1[7] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3448 = io_in_bits_DecodeIn_data_src1[8] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3450 = io_in_bits_DecodeIn_data_src1[9] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3452 = io_in_bits_DecodeIn_data_src1[10] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3454 = io_in_bits_DecodeIn_data_src1[11] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3456 = io_in_bits_DecodeIn_data_src1[12] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3458 = io_in_bits_DecodeIn_data_src1[13] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3460 = io_in_bits_DecodeIn_data_src1[14] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3462 = io_in_bits_DecodeIn_data_src1[15] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3464 = io_in_bits_DecodeIn_data_src1[16] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3466 = io_in_bits_DecodeIn_data_src1[17] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3468 = io_in_bits_DecodeIn_data_src1[18] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3470 = io_in_bits_DecodeIn_data_src1[19] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3472 = io_in_bits_DecodeIn_data_src1[20] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3474 = io_in_bits_DecodeIn_data_src1[21] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3476 = io_in_bits_DecodeIn_data_src1[22] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3478 = io_in_bits_DecodeIn_data_src1[23] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3480 = io_in_bits_DecodeIn_data_src1[24] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3482 = io_in_bits_DecodeIn_data_src1[25] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3484 = io_in_bits_DecodeIn_data_src1[26] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3486 = io_in_bits_DecodeIn_data_src1[27] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3488 = io_in_bits_DecodeIn_data_src1[28] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3490 = io_in_bits_DecodeIn_data_src1[29] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3492 = io_in_bits_DecodeIn_data_src1[30] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3494 = io_in_bits_DecodeIn_data_src1[31] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3496 = _T_3492 & _T_3494; // @[PALU.scala 427:113]
  wire  _T_3498 = _T_3490 & (_T_3492 & _T_3494); // @[PALU.scala 427:113]
  wire  _T_3500 = _T_3488 & (_T_3490 & (_T_3492 & _T_3494)); // @[PALU.scala 427:113]
  wire  _T_3502 = _T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))); // @[PALU.scala 427:113]
  wire  _T_3504 = _T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))); // @[PALU.scala 427:113]
  wire  _T_3506 = _T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))); // @[PALU.scala 427:113]
  wire  _T_3508 = _T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))); // @[PALU.scala 427:113]
  wire  _T_3510 = _T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))); // @[PALU.scala 427:113]
  wire  _T_3512 = _T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 &
    _T_3494)))))))); // @[PALU.scala 427:113]
  wire  _T_3514 = _T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (
    _T_3492 & _T_3494))))))))); // @[PALU.scala 427:113]
  wire  _T_3516 = _T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (
    _T_3490 & (_T_3492 & _T_3494)))))))))); // @[PALU.scala 427:113]
  wire  _T_3518 = _T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (
    _T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))); // @[PALU.scala 427:113]
  wire  _T_3520 = _T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (
    _T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))); // @[PALU.scala 427:113]
  wire  _T_3522 = _T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (
    _T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3524 = _T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (
    _T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3526 = _T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (
    _T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3528 = _T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (
    _T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3530 = _T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (
    _T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))
    )))))); // @[PALU.scala 427:113]
  wire  _T_3532 = _T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (
    _T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494
    )))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3534 = _T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (
    _T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (
    _T_3492 & _T_3494))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3536 = _T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (
    _T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (
    _T_3490 & (_T_3492 & _T_3494)))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3538 = _T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (
    _T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (
    _T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3540 = _T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (
    _T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (
    _T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3542 = _T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (
    _T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (
    _T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3544 = _T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (
    _T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (
    _T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3546 = _T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (
    _T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (
    _T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3548 = _T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (
    _T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (
    _T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))))
    )))); // @[PALU.scala 427:113]
  wire  _T_3550 = _T_3438 & (_T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (
    _T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (
    _T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))
    )))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3552 = _T_3436 & (_T_3438 & (_T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (
    _T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (
    _T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494
    )))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3554 = _T_3434 & (_T_3436 & (_T_3438 & (_T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (
    _T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (
    _T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (
    _T_3492 & _T_3494))))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3556 = _T_3432 & _T_3554; // @[PALU.scala 427:113]
  wire [1:0] _T_3557 = _T_3494 + _T_3496; // @[PALU.scala 428:38]
  wire [1:0] _GEN_759 = {{1'd0}, _T_3498}; // @[PALU.scala 428:38]
  wire [2:0] _T_3558 = _T_3557 + _GEN_759; // @[PALU.scala 428:38]
  wire [2:0] _GEN_760 = {{2'd0}, _T_3500}; // @[PALU.scala 428:38]
  wire [3:0] _T_3559 = _T_3558 + _GEN_760; // @[PALU.scala 428:38]
  wire [3:0] _GEN_761 = {{3'd0}, _T_3502}; // @[PALU.scala 428:38]
  wire [4:0] _T_3560 = _T_3559 + _GEN_761; // @[PALU.scala 428:38]
  wire [4:0] _GEN_762 = {{4'd0}, _T_3504}; // @[PALU.scala 428:38]
  wire [5:0] _T_3561 = _T_3560 + _GEN_762; // @[PALU.scala 428:38]
  wire [5:0] _GEN_763 = {{5'd0}, _T_3506}; // @[PALU.scala 428:38]
  wire [6:0] _T_3562 = _T_3561 + _GEN_763; // @[PALU.scala 428:38]
  wire [6:0] _GEN_764 = {{6'd0}, _T_3508}; // @[PALU.scala 428:38]
  wire [7:0] _T_3563 = _T_3562 + _GEN_764; // @[PALU.scala 428:38]
  wire [7:0] _GEN_765 = {{7'd0}, _T_3510}; // @[PALU.scala 428:38]
  wire [8:0] _T_3564 = _T_3563 + _GEN_765; // @[PALU.scala 428:38]
  wire [8:0] _GEN_766 = {{8'd0}, _T_3512}; // @[PALU.scala 428:38]
  wire [9:0] _T_3565 = _T_3564 + _GEN_766; // @[PALU.scala 428:38]
  wire [9:0] _GEN_767 = {{9'd0}, _T_3514}; // @[PALU.scala 428:38]
  wire [10:0] _T_3566 = _T_3565 + _GEN_767; // @[PALU.scala 428:38]
  wire [10:0] _GEN_768 = {{10'd0}, _T_3516}; // @[PALU.scala 428:38]
  wire [11:0] _T_3567 = _T_3566 + _GEN_768; // @[PALU.scala 428:38]
  wire [11:0] _GEN_769 = {{11'd0}, _T_3518}; // @[PALU.scala 428:38]
  wire [12:0] _T_3568 = _T_3567 + _GEN_769; // @[PALU.scala 428:38]
  wire [12:0] _GEN_770 = {{12'd0}, _T_3520}; // @[PALU.scala 428:38]
  wire [13:0] _T_3569 = _T_3568 + _GEN_770; // @[PALU.scala 428:38]
  wire [13:0] _GEN_771 = {{13'd0}, _T_3522}; // @[PALU.scala 428:38]
  wire [14:0] _T_3570 = _T_3569 + _GEN_771; // @[PALU.scala 428:38]
  wire [14:0] _GEN_772 = {{14'd0}, _T_3524}; // @[PALU.scala 428:38]
  wire [15:0] _T_3571 = _T_3570 + _GEN_772; // @[PALU.scala 428:38]
  wire [15:0] _GEN_773 = {{15'd0}, _T_3526}; // @[PALU.scala 428:38]
  wire [16:0] _T_3572 = _T_3571 + _GEN_773; // @[PALU.scala 428:38]
  wire [16:0] _GEN_774 = {{16'd0}, _T_3528}; // @[PALU.scala 428:38]
  wire [17:0] _T_3573 = _T_3572 + _GEN_774; // @[PALU.scala 428:38]
  wire [17:0] _GEN_775 = {{17'd0}, _T_3530}; // @[PALU.scala 428:38]
  wire [18:0] _T_3574 = _T_3573 + _GEN_775; // @[PALU.scala 428:38]
  wire [18:0] _GEN_776 = {{18'd0}, _T_3532}; // @[PALU.scala 428:38]
  wire [19:0] _T_3575 = _T_3574 + _GEN_776; // @[PALU.scala 428:38]
  wire [19:0] _GEN_777 = {{19'd0}, _T_3534}; // @[PALU.scala 428:38]
  wire [20:0] _T_3576 = _T_3575 + _GEN_777; // @[PALU.scala 428:38]
  wire [20:0] _GEN_778 = {{20'd0}, _T_3536}; // @[PALU.scala 428:38]
  wire [21:0] _T_3577 = _T_3576 + _GEN_778; // @[PALU.scala 428:38]
  wire [21:0] _GEN_779 = {{21'd0}, _T_3538}; // @[PALU.scala 428:38]
  wire [22:0] _T_3578 = _T_3577 + _GEN_779; // @[PALU.scala 428:38]
  wire [22:0] _GEN_780 = {{22'd0}, _T_3540}; // @[PALU.scala 428:38]
  wire [23:0] _T_3579 = _T_3578 + _GEN_780; // @[PALU.scala 428:38]
  wire [23:0] _GEN_781 = {{23'd0}, _T_3542}; // @[PALU.scala 428:38]
  wire [24:0] _T_3580 = _T_3579 + _GEN_781; // @[PALU.scala 428:38]
  wire [24:0] _GEN_782 = {{24'd0}, _T_3544}; // @[PALU.scala 428:38]
  wire [25:0] _T_3581 = _T_3580 + _GEN_782; // @[PALU.scala 428:38]
  wire [25:0] _GEN_783 = {{25'd0}, _T_3546}; // @[PALU.scala 428:38]
  wire [26:0] _T_3582 = _T_3581 + _GEN_783; // @[PALU.scala 428:38]
  wire [26:0] _GEN_784 = {{26'd0}, _T_3548}; // @[PALU.scala 428:38]
  wire [27:0] _T_3583 = _T_3582 + _GEN_784; // @[PALU.scala 428:38]
  wire [27:0] _GEN_785 = {{27'd0}, _T_3550}; // @[PALU.scala 428:38]
  wire [28:0] _T_3584 = _T_3583 + _GEN_785; // @[PALU.scala 428:38]
  wire [28:0] _GEN_786 = {{28'd0}, _T_3552}; // @[PALU.scala 428:38]
  wire [29:0] _T_3585 = _T_3584 + _GEN_786; // @[PALU.scala 428:38]
  wire [29:0] _GEN_787 = {{29'd0}, _T_3554}; // @[PALU.scala 428:38]
  wire [30:0] _T_3586 = _T_3585 + _GEN_787; // @[PALU.scala 428:38]
  wire [30:0] _GEN_788 = {{30'd0}, _T_3556}; // @[PALU.scala 428:38]
  wire [31:0] _T_3587 = _T_3586 + _GEN_788; // @[PALU.scala 428:38]
  wire [31:0] _T_3589 = _T_3587 - 32'h1; // @[PALU.scala 429:44]
  wire [31:0] _T_3590 = io_in_bits_DecodeIn_data_src2[0] ? _T_3587 : _T_3589; // @[PALU.scala 429:26]
  wire  _T_3593 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[63]; // @[PALU.scala 423:29]
  wire  _T_3595 = io_in_bits_DecodeIn_data_src1[32] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3597 = io_in_bits_DecodeIn_data_src1[33] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3599 = io_in_bits_DecodeIn_data_src1[34] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3601 = io_in_bits_DecodeIn_data_src1[35] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3603 = io_in_bits_DecodeIn_data_src1[36] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3605 = io_in_bits_DecodeIn_data_src1[37] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3607 = io_in_bits_DecodeIn_data_src1[38] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3609 = io_in_bits_DecodeIn_data_src1[39] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3611 = io_in_bits_DecodeIn_data_src1[40] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3613 = io_in_bits_DecodeIn_data_src1[41] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3615 = io_in_bits_DecodeIn_data_src1[42] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3617 = io_in_bits_DecodeIn_data_src1[43] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3619 = io_in_bits_DecodeIn_data_src1[44] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3621 = io_in_bits_DecodeIn_data_src1[45] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3623 = io_in_bits_DecodeIn_data_src1[46] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3625 = io_in_bits_DecodeIn_data_src1[47] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3627 = io_in_bits_DecodeIn_data_src1[48] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3629 = io_in_bits_DecodeIn_data_src1[49] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3631 = io_in_bits_DecodeIn_data_src1[50] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3633 = io_in_bits_DecodeIn_data_src1[51] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3635 = io_in_bits_DecodeIn_data_src1[52] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3637 = io_in_bits_DecodeIn_data_src1[53] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3639 = io_in_bits_DecodeIn_data_src1[54] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3641 = io_in_bits_DecodeIn_data_src1[55] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3643 = io_in_bits_DecodeIn_data_src1[56] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3645 = io_in_bits_DecodeIn_data_src1[57] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3647 = io_in_bits_DecodeIn_data_src1[58] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3649 = io_in_bits_DecodeIn_data_src1[59] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3651 = io_in_bits_DecodeIn_data_src1[60] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3653 = io_in_bits_DecodeIn_data_src1[61] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3655 = io_in_bits_DecodeIn_data_src1[62] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3657 = io_in_bits_DecodeIn_data_src1[63] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3659 = _T_3655 & _T_3657; // @[PALU.scala 427:113]
  wire  _T_3661 = _T_3653 & (_T_3655 & _T_3657); // @[PALU.scala 427:113]
  wire  _T_3663 = _T_3651 & (_T_3653 & (_T_3655 & _T_3657)); // @[PALU.scala 427:113]
  wire  _T_3665 = _T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))); // @[PALU.scala 427:113]
  wire  _T_3667 = _T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))); // @[PALU.scala 427:113]
  wire  _T_3669 = _T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))); // @[PALU.scala 427:113]
  wire  _T_3671 = _T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))); // @[PALU.scala 427:113]
  wire  _T_3673 = _T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))); // @[PALU.scala 427:113]
  wire  _T_3675 = _T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 &
    _T_3657)))))))); // @[PALU.scala 427:113]
  wire  _T_3677 = _T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (
    _T_3655 & _T_3657))))))))); // @[PALU.scala 427:113]
  wire  _T_3679 = _T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (
    _T_3653 & (_T_3655 & _T_3657)))))))))); // @[PALU.scala 427:113]
  wire  _T_3681 = _T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (
    _T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))); // @[PALU.scala 427:113]
  wire  _T_3683 = _T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (
    _T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))); // @[PALU.scala 427:113]
  wire  _T_3685 = _T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (
    _T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3687 = _T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (
    _T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3689 = _T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (
    _T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3691 = _T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (
    _T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3693 = _T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (
    _T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))
    )))))); // @[PALU.scala 427:113]
  wire  _T_3695 = _T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (
    _T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657
    )))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3697 = _T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (
    _T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (
    _T_3655 & _T_3657))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3699 = _T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (
    _T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (
    _T_3653 & (_T_3655 & _T_3657)))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3701 = _T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (
    _T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (
    _T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3703 = _T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (
    _T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (
    _T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3705 = _T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (
    _T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (
    _T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3707 = _T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (
    _T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (
    _T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3709 = _T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (
    _T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (
    _T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3711 = _T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (
    _T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (
    _T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))))
    )))); // @[PALU.scala 427:113]
  wire  _T_3713 = _T_3601 & (_T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (
    _T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (
    _T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))
    )))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3715 = _T_3599 & (_T_3601 & (_T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (
    _T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (
    _T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657
    )))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3717 = _T_3597 & (_T_3599 & (_T_3601 & (_T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (
    _T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (
    _T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (
    _T_3655 & _T_3657))))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3719 = _T_3595 & _T_3717; // @[PALU.scala 427:113]
  wire [1:0] _T_3720 = _T_3657 + _T_3659; // @[PALU.scala 428:38]
  wire [1:0] _GEN_789 = {{1'd0}, _T_3661}; // @[PALU.scala 428:38]
  wire [2:0] _T_3721 = _T_3720 + _GEN_789; // @[PALU.scala 428:38]
  wire [2:0] _GEN_790 = {{2'd0}, _T_3663}; // @[PALU.scala 428:38]
  wire [3:0] _T_3722 = _T_3721 + _GEN_790; // @[PALU.scala 428:38]
  wire [3:0] _GEN_791 = {{3'd0}, _T_3665}; // @[PALU.scala 428:38]
  wire [4:0] _T_3723 = _T_3722 + _GEN_791; // @[PALU.scala 428:38]
  wire [4:0] _GEN_792 = {{4'd0}, _T_3667}; // @[PALU.scala 428:38]
  wire [5:0] _T_3724 = _T_3723 + _GEN_792; // @[PALU.scala 428:38]
  wire [5:0] _GEN_793 = {{5'd0}, _T_3669}; // @[PALU.scala 428:38]
  wire [6:0] _T_3725 = _T_3724 + _GEN_793; // @[PALU.scala 428:38]
  wire [6:0] _GEN_794 = {{6'd0}, _T_3671}; // @[PALU.scala 428:38]
  wire [7:0] _T_3726 = _T_3725 + _GEN_794; // @[PALU.scala 428:38]
  wire [7:0] _GEN_795 = {{7'd0}, _T_3673}; // @[PALU.scala 428:38]
  wire [8:0] _T_3727 = _T_3726 + _GEN_795; // @[PALU.scala 428:38]
  wire [8:0] _GEN_796 = {{8'd0}, _T_3675}; // @[PALU.scala 428:38]
  wire [9:0] _T_3728 = _T_3727 + _GEN_796; // @[PALU.scala 428:38]
  wire [9:0] _GEN_797 = {{9'd0}, _T_3677}; // @[PALU.scala 428:38]
  wire [10:0] _T_3729 = _T_3728 + _GEN_797; // @[PALU.scala 428:38]
  wire [10:0] _GEN_798 = {{10'd0}, _T_3679}; // @[PALU.scala 428:38]
  wire [11:0] _T_3730 = _T_3729 + _GEN_798; // @[PALU.scala 428:38]
  wire [11:0] _GEN_799 = {{11'd0}, _T_3681}; // @[PALU.scala 428:38]
  wire [12:0] _T_3731 = _T_3730 + _GEN_799; // @[PALU.scala 428:38]
  wire [12:0] _GEN_800 = {{12'd0}, _T_3683}; // @[PALU.scala 428:38]
  wire [13:0] _T_3732 = _T_3731 + _GEN_800; // @[PALU.scala 428:38]
  wire [13:0] _GEN_801 = {{13'd0}, _T_3685}; // @[PALU.scala 428:38]
  wire [14:0] _T_3733 = _T_3732 + _GEN_801; // @[PALU.scala 428:38]
  wire [14:0] _GEN_802 = {{14'd0}, _T_3687}; // @[PALU.scala 428:38]
  wire [15:0] _T_3734 = _T_3733 + _GEN_802; // @[PALU.scala 428:38]
  wire [15:0] _GEN_803 = {{15'd0}, _T_3689}; // @[PALU.scala 428:38]
  wire [16:0] _T_3735 = _T_3734 + _GEN_803; // @[PALU.scala 428:38]
  wire [16:0] _GEN_804 = {{16'd0}, _T_3691}; // @[PALU.scala 428:38]
  wire [17:0] _T_3736 = _T_3735 + _GEN_804; // @[PALU.scala 428:38]
  wire [17:0] _GEN_805 = {{17'd0}, _T_3693}; // @[PALU.scala 428:38]
  wire [18:0] _T_3737 = _T_3736 + _GEN_805; // @[PALU.scala 428:38]
  wire [18:0] _GEN_806 = {{18'd0}, _T_3695}; // @[PALU.scala 428:38]
  wire [19:0] _T_3738 = _T_3737 + _GEN_806; // @[PALU.scala 428:38]
  wire [19:0] _GEN_807 = {{19'd0}, _T_3697}; // @[PALU.scala 428:38]
  wire [20:0] _T_3739 = _T_3738 + _GEN_807; // @[PALU.scala 428:38]
  wire [20:0] _GEN_808 = {{20'd0}, _T_3699}; // @[PALU.scala 428:38]
  wire [21:0] _T_3740 = _T_3739 + _GEN_808; // @[PALU.scala 428:38]
  wire [21:0] _GEN_809 = {{21'd0}, _T_3701}; // @[PALU.scala 428:38]
  wire [22:0] _T_3741 = _T_3740 + _GEN_809; // @[PALU.scala 428:38]
  wire [22:0] _GEN_810 = {{22'd0}, _T_3703}; // @[PALU.scala 428:38]
  wire [23:0] _T_3742 = _T_3741 + _GEN_810; // @[PALU.scala 428:38]
  wire [23:0] _GEN_811 = {{23'd0}, _T_3705}; // @[PALU.scala 428:38]
  wire [24:0] _T_3743 = _T_3742 + _GEN_811; // @[PALU.scala 428:38]
  wire [24:0] _GEN_812 = {{24'd0}, _T_3707}; // @[PALU.scala 428:38]
  wire [25:0] _T_3744 = _T_3743 + _GEN_812; // @[PALU.scala 428:38]
  wire [25:0] _GEN_813 = {{25'd0}, _T_3709}; // @[PALU.scala 428:38]
  wire [26:0] _T_3745 = _T_3744 + _GEN_813; // @[PALU.scala 428:38]
  wire [26:0] _GEN_814 = {{26'd0}, _T_3711}; // @[PALU.scala 428:38]
  wire [27:0] _T_3746 = _T_3745 + _GEN_814; // @[PALU.scala 428:38]
  wire [27:0] _GEN_815 = {{27'd0}, _T_3713}; // @[PALU.scala 428:38]
  wire [28:0] _T_3747 = _T_3746 + _GEN_815; // @[PALU.scala 428:38]
  wire [28:0] _GEN_816 = {{28'd0}, _T_3715}; // @[PALU.scala 428:38]
  wire [29:0] _T_3748 = _T_3747 + _GEN_816; // @[PALU.scala 428:38]
  wire [29:0] _GEN_817 = {{29'd0}, _T_3717}; // @[PALU.scala 428:38]
  wire [30:0] _T_3749 = _T_3748 + _GEN_817; // @[PALU.scala 428:38]
  wire [30:0] _GEN_818 = {{30'd0}, _T_3719}; // @[PALU.scala 428:38]
  wire [31:0] _T_3750 = _T_3749 + _GEN_818; // @[PALU.scala 428:38]
  wire [31:0] _T_3752 = _T_3750 - 32'h1; // @[PALU.scala 429:44]
  wire [31:0] _T_3753 = io_in_bits_DecodeIn_data_src2[0] ? _T_3750 : _T_3752; // @[PALU.scala 429:26]
  wire [63:0] _T_3754 = {_T_3753,_T_3590}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_555 = io_in_bits_Pctrl_isCnt_32 ? _T_3754 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 577:25 579:16]
  wire [63:0] _GEN_556 = io_in_bits_Pctrl_isCnt_8 ? _T_3425 : _GEN_555; // @[PALU.scala 574:24 576:16]
  wire [63:0] cntRes = io_in_bits_Pctrl_isCnt_16 ? _T_3072 : _GEN_556; // @[PALU.scala 571:19 573:16]
  wire [15:0] _GEN_558 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src1[31:16] : 16'h0; // @[PALU.scala 450:37 451:24]
  wire [15:0] _GEN_559 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src2[31:16] : 16'h0; // @[PALU.scala 450:37 452:24]
  wire [15:0] _GEN_560 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src1[31:16] :
    _GEN_558; // @[PALU.scala 447:37 448:24]
  wire [15:0] _GEN_561 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src2[15:0] : _GEN_559
    ; // @[PALU.scala 447:37 449:24]
  wire [15:0] _GEN_562 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src1[15:0] : _GEN_560
    ; // @[PALU.scala 443:37 444:24]
  wire [15:0] _GEN_563 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src2[31:16] :
    _GEN_561; // @[PALU.scala 443:37 445:24]
  wire [15:0] _GEN_564 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src1[15:0] : _GEN_562
    ; // @[PALU.scala 440:31 441:24]
  wire [15:0] _GEN_565 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src2[15:0] : _GEN_563
    ; // @[PALU.scala 440:31 442:24]
  wire [15:0] _GEN_566 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src1[63:48] : 16'h0; // @[PALU.scala 450:37 451:24]
  wire [15:0] _GEN_567 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src2[63:48] : 16'h0; // @[PALU.scala 450:37 452:24]
  wire [15:0] _GEN_568 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src1[63:48] :
    _GEN_566; // @[PALU.scala 447:37 448:24]
  wire [15:0] _GEN_569 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src2[47:32] :
    _GEN_567; // @[PALU.scala 447:37 449:24]
  wire [15:0] _GEN_570 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src1[47:32] :
    _GEN_568; // @[PALU.scala 443:37 444:24]
  wire [15:0] _GEN_571 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src2[63:48] :
    _GEN_569; // @[PALU.scala 443:37 445:24]
  wire [15:0] _GEN_572 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src1[47:32] :
    _GEN_570; // @[PALU.scala 440:31 441:24]
  wire [15:0] _GEN_573 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src2[47:32] :
    _GEN_571; // @[PALU.scala 440:31 442:24]
  wire [63:0] _T_3841 = {_GEN_572,_GEN_573,_GEN_564,_GEN_565}; // @[Cat.scala 30:58]
  wire [63:0] _T_4012 = {io_in_bits_DecodeIn_data_src1[55:48],io_in_bits_DecodeIn_data_src1[63:56],
    io_in_bits_DecodeIn_data_src1[39:32],io_in_bits_DecodeIn_data_src1[47:40],io_in_bits_DecodeIn_data_src1[23:16],
    io_in_bits_DecodeIn_data_src1[31:24],io_in_bits_DecodeIn_data_src1[7:0],io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_606 = io_in_bits_Pctrl_isSwap_8 ? _T_4012 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 586:25 587:17]
  wire [63:0] swapRes = io_in_bits_Pctrl_isSwap_16 ? _T_3841 : _GEN_606; // @[PALU.scala 584:20 585:17]
  wire [63:0] _GEN_819 = {{32'd0}, io_in_bits_DecodeIn_data_src1[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4016 = _GEN_819 & 64'hffffffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4018 = {io_in_bits_DecodeIn_data_src1[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4020 = _T_4018 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4021 = _T_4016 | _T_4020; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_820 = {{16'd0}, _T_4021[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4026 = _GEN_820 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4028 = {_T_4021[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4030 = _T_4028 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4031 = _T_4026 | _T_4030; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_821 = {{8'd0}, _T_4031[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4036 = _GEN_821 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4038 = {_T_4031[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4040 = _T_4038 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4041 = _T_4036 | _T_4040; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_822 = {{4'd0}, _T_4041[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4046 = _GEN_822 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4048 = {_T_4041[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4050 = _T_4048 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4051 = _T_4046 | _T_4050; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_823 = {{2'd0}, _T_4051[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4056 = _GEN_823 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4058 = {_T_4051[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4060 = _T_4058 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4061 = _T_4056 | _T_4060; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_824 = {{1'd0}, _T_4061[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4066 = _GEN_824 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4068 = {_T_4061[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4070 = _T_4068 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4071 = _T_4066 | _T_4070; // @[Bitwise.scala 103:39]
  wire [63:0] bitrevRes = io_in_bits_Pctrl_isBitrev ? _T_4071 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 592:19 593:19]
  wire  _T_4077 = io_in_bits_DecodeIn_data_src2[0] ? io_in_bits_DecodeIn_data_src1[0] : io_in_bits_DecodeIn_data_src3[0]
    ; // @[PALU.scala 477:46]
  wire  _T_4082 = io_in_bits_DecodeIn_data_src2[1] ? io_in_bits_DecodeIn_data_src1[1] : io_in_bits_DecodeIn_data_src3[1]
    ; // @[PALU.scala 477:46]
  wire  _T_4087 = io_in_bits_DecodeIn_data_src2[2] ? io_in_bits_DecodeIn_data_src1[2] : io_in_bits_DecodeIn_data_src3[2]
    ; // @[PALU.scala 477:46]
  wire  _T_4092 = io_in_bits_DecodeIn_data_src2[3] ? io_in_bits_DecodeIn_data_src1[3] : io_in_bits_DecodeIn_data_src3[3]
    ; // @[PALU.scala 477:46]
  wire  _T_4097 = io_in_bits_DecodeIn_data_src2[4] ? io_in_bits_DecodeIn_data_src1[4] : io_in_bits_DecodeIn_data_src3[4]
    ; // @[PALU.scala 477:46]
  wire  _T_4102 = io_in_bits_DecodeIn_data_src2[5] ? io_in_bits_DecodeIn_data_src1[5] : io_in_bits_DecodeIn_data_src3[5]
    ; // @[PALU.scala 477:46]
  wire  _T_4107 = io_in_bits_DecodeIn_data_src2[6] ? io_in_bits_DecodeIn_data_src1[6] : io_in_bits_DecodeIn_data_src3[6]
    ; // @[PALU.scala 477:46]
  wire  _T_4112 = io_in_bits_DecodeIn_data_src2[7] ? io_in_bits_DecodeIn_data_src1[7] : io_in_bits_DecodeIn_data_src3[7]
    ; // @[PALU.scala 477:46]
  wire  _T_4117 = io_in_bits_DecodeIn_data_src2[8] ? io_in_bits_DecodeIn_data_src1[8] : io_in_bits_DecodeIn_data_src3[8]
    ; // @[PALU.scala 477:46]
  wire  _T_4122 = io_in_bits_DecodeIn_data_src2[9] ? io_in_bits_DecodeIn_data_src1[9] : io_in_bits_DecodeIn_data_src3[9]
    ; // @[PALU.scala 477:46]
  wire  _T_4127 = io_in_bits_DecodeIn_data_src2[10] ? io_in_bits_DecodeIn_data_src1[10] : io_in_bits_DecodeIn_data_src3[
    10]; // @[PALU.scala 477:46]
  wire  _T_4132 = io_in_bits_DecodeIn_data_src2[11] ? io_in_bits_DecodeIn_data_src1[11] : io_in_bits_DecodeIn_data_src3[
    11]; // @[PALU.scala 477:46]
  wire  _T_4137 = io_in_bits_DecodeIn_data_src2[12] ? io_in_bits_DecodeIn_data_src1[12] : io_in_bits_DecodeIn_data_src3[
    12]; // @[PALU.scala 477:46]
  wire  _T_4142 = io_in_bits_DecodeIn_data_src2[13] ? io_in_bits_DecodeIn_data_src1[13] : io_in_bits_DecodeIn_data_src3[
    13]; // @[PALU.scala 477:46]
  wire  _T_4147 = io_in_bits_DecodeIn_data_src2[14] ? io_in_bits_DecodeIn_data_src1[14] : io_in_bits_DecodeIn_data_src3[
    14]; // @[PALU.scala 477:46]
  wire  _T_4152 = io_in_bits_DecodeIn_data_src2[15] ? io_in_bits_DecodeIn_data_src1[15] : io_in_bits_DecodeIn_data_src3[
    15]; // @[PALU.scala 477:46]
  wire  _T_4157 = io_in_bits_DecodeIn_data_src2[16] ? io_in_bits_DecodeIn_data_src1[16] : io_in_bits_DecodeIn_data_src3[
    16]; // @[PALU.scala 477:46]
  wire  _T_4162 = io_in_bits_DecodeIn_data_src2[17] ? io_in_bits_DecodeIn_data_src1[17] : io_in_bits_DecodeIn_data_src3[
    17]; // @[PALU.scala 477:46]
  wire  _T_4167 = io_in_bits_DecodeIn_data_src2[18] ? io_in_bits_DecodeIn_data_src1[18] : io_in_bits_DecodeIn_data_src3[
    18]; // @[PALU.scala 477:46]
  wire  _T_4172 = io_in_bits_DecodeIn_data_src2[19] ? io_in_bits_DecodeIn_data_src1[19] : io_in_bits_DecodeIn_data_src3[
    19]; // @[PALU.scala 477:46]
  wire  _T_4177 = io_in_bits_DecodeIn_data_src2[20] ? io_in_bits_DecodeIn_data_src1[20] : io_in_bits_DecodeIn_data_src3[
    20]; // @[PALU.scala 477:46]
  wire  _T_4182 = io_in_bits_DecodeIn_data_src2[21] ? io_in_bits_DecodeIn_data_src1[21] : io_in_bits_DecodeIn_data_src3[
    21]; // @[PALU.scala 477:46]
  wire  _T_4187 = io_in_bits_DecodeIn_data_src2[22] ? io_in_bits_DecodeIn_data_src1[22] : io_in_bits_DecodeIn_data_src3[
    22]; // @[PALU.scala 477:46]
  wire  _T_4192 = io_in_bits_DecodeIn_data_src2[23] ? io_in_bits_DecodeIn_data_src1[23] : io_in_bits_DecodeIn_data_src3[
    23]; // @[PALU.scala 477:46]
  wire  _T_4197 = io_in_bits_DecodeIn_data_src2[24] ? io_in_bits_DecodeIn_data_src1[24] : io_in_bits_DecodeIn_data_src3[
    24]; // @[PALU.scala 477:46]
  wire  _T_4202 = io_in_bits_DecodeIn_data_src2[25] ? io_in_bits_DecodeIn_data_src1[25] : io_in_bits_DecodeIn_data_src3[
    25]; // @[PALU.scala 477:46]
  wire  _T_4207 = io_in_bits_DecodeIn_data_src2[26] ? io_in_bits_DecodeIn_data_src1[26] : io_in_bits_DecodeIn_data_src3[
    26]; // @[PALU.scala 477:46]
  wire  _T_4212 = io_in_bits_DecodeIn_data_src2[27] ? io_in_bits_DecodeIn_data_src1[27] : io_in_bits_DecodeIn_data_src3[
    27]; // @[PALU.scala 477:46]
  wire  _T_4217 = io_in_bits_DecodeIn_data_src2[28] ? io_in_bits_DecodeIn_data_src1[28] : io_in_bits_DecodeIn_data_src3[
    28]; // @[PALU.scala 477:46]
  wire  _T_4222 = io_in_bits_DecodeIn_data_src2[29] ? io_in_bits_DecodeIn_data_src1[29] : io_in_bits_DecodeIn_data_src3[
    29]; // @[PALU.scala 477:46]
  wire  _T_4227 = io_in_bits_DecodeIn_data_src2[30] ? io_in_bits_DecodeIn_data_src1[30] : io_in_bits_DecodeIn_data_src3[
    30]; // @[PALU.scala 477:46]
  wire  _T_4232 = io_in_bits_DecodeIn_data_src2[31] ? io_in_bits_DecodeIn_data_src1[31] : io_in_bits_DecodeIn_data_src3[
    31]; // @[PALU.scala 477:46]
  wire  _T_4237 = io_in_bits_DecodeIn_data_src2[32] ? io_in_bits_DecodeIn_data_src1[32] : io_in_bits_DecodeIn_data_src3[
    32]; // @[PALU.scala 477:46]
  wire  _T_4242 = io_in_bits_DecodeIn_data_src2[33] ? io_in_bits_DecodeIn_data_src1[33] : io_in_bits_DecodeIn_data_src3[
    33]; // @[PALU.scala 477:46]
  wire  _T_4247 = io_in_bits_DecodeIn_data_src2[34] ? io_in_bits_DecodeIn_data_src1[34] : io_in_bits_DecodeIn_data_src3[
    34]; // @[PALU.scala 477:46]
  wire  _T_4252 = io_in_bits_DecodeIn_data_src2[35] ? io_in_bits_DecodeIn_data_src1[35] : io_in_bits_DecodeIn_data_src3[
    35]; // @[PALU.scala 477:46]
  wire  _T_4257 = io_in_bits_DecodeIn_data_src2[36] ? io_in_bits_DecodeIn_data_src1[36] : io_in_bits_DecodeIn_data_src3[
    36]; // @[PALU.scala 477:46]
  wire  _T_4262 = io_in_bits_DecodeIn_data_src2[37] ? io_in_bits_DecodeIn_data_src1[37] : io_in_bits_DecodeIn_data_src3[
    37]; // @[PALU.scala 477:46]
  wire  _T_4267 = io_in_bits_DecodeIn_data_src2[38] ? io_in_bits_DecodeIn_data_src1[38] : io_in_bits_DecodeIn_data_src3[
    38]; // @[PALU.scala 477:46]
  wire  _T_4272 = io_in_bits_DecodeIn_data_src2[39] ? io_in_bits_DecodeIn_data_src1[39] : io_in_bits_DecodeIn_data_src3[
    39]; // @[PALU.scala 477:46]
  wire  _T_4277 = io_in_bits_DecodeIn_data_src2[40] ? io_in_bits_DecodeIn_data_src1[40] : io_in_bits_DecodeIn_data_src3[
    40]; // @[PALU.scala 477:46]
  wire  _T_4282 = io_in_bits_DecodeIn_data_src2[41] ? io_in_bits_DecodeIn_data_src1[41] : io_in_bits_DecodeIn_data_src3[
    41]; // @[PALU.scala 477:46]
  wire  _T_4287 = io_in_bits_DecodeIn_data_src2[42] ? io_in_bits_DecodeIn_data_src1[42] : io_in_bits_DecodeIn_data_src3[
    42]; // @[PALU.scala 477:46]
  wire  _T_4292 = io_in_bits_DecodeIn_data_src2[43] ? io_in_bits_DecodeIn_data_src1[43] : io_in_bits_DecodeIn_data_src3[
    43]; // @[PALU.scala 477:46]
  wire  _T_4297 = io_in_bits_DecodeIn_data_src2[44] ? io_in_bits_DecodeIn_data_src1[44] : io_in_bits_DecodeIn_data_src3[
    44]; // @[PALU.scala 477:46]
  wire  _T_4302 = io_in_bits_DecodeIn_data_src2[45] ? io_in_bits_DecodeIn_data_src1[45] : io_in_bits_DecodeIn_data_src3[
    45]; // @[PALU.scala 477:46]
  wire  _T_4307 = io_in_bits_DecodeIn_data_src2[46] ? io_in_bits_DecodeIn_data_src1[46] : io_in_bits_DecodeIn_data_src3[
    46]; // @[PALU.scala 477:46]
  wire  _T_4312 = io_in_bits_DecodeIn_data_src2[47] ? io_in_bits_DecodeIn_data_src1[47] : io_in_bits_DecodeIn_data_src3[
    47]; // @[PALU.scala 477:46]
  wire  _T_4317 = io_in_bits_DecodeIn_data_src2[48] ? io_in_bits_DecodeIn_data_src1[48] : io_in_bits_DecodeIn_data_src3[
    48]; // @[PALU.scala 477:46]
  wire  _T_4322 = io_in_bits_DecodeIn_data_src2[49] ? io_in_bits_DecodeIn_data_src1[49] : io_in_bits_DecodeIn_data_src3[
    49]; // @[PALU.scala 477:46]
  wire  _T_4327 = io_in_bits_DecodeIn_data_src2[50] ? io_in_bits_DecodeIn_data_src1[50] : io_in_bits_DecodeIn_data_src3[
    50]; // @[PALU.scala 477:46]
  wire  _T_4332 = io_in_bits_DecodeIn_data_src2[51] ? io_in_bits_DecodeIn_data_src1[51] : io_in_bits_DecodeIn_data_src3[
    51]; // @[PALU.scala 477:46]
  wire  _T_4337 = io_in_bits_DecodeIn_data_src2[52] ? io_in_bits_DecodeIn_data_src1[52] : io_in_bits_DecodeIn_data_src3[
    52]; // @[PALU.scala 477:46]
  wire  _T_4342 = io_in_bits_DecodeIn_data_src2[53] ? io_in_bits_DecodeIn_data_src1[53] : io_in_bits_DecodeIn_data_src3[
    53]; // @[PALU.scala 477:46]
  wire  _T_4347 = io_in_bits_DecodeIn_data_src2[54] ? io_in_bits_DecodeIn_data_src1[54] : io_in_bits_DecodeIn_data_src3[
    54]; // @[PALU.scala 477:46]
  wire  _T_4352 = io_in_bits_DecodeIn_data_src2[55] ? io_in_bits_DecodeIn_data_src1[55] : io_in_bits_DecodeIn_data_src3[
    55]; // @[PALU.scala 477:46]
  wire  _T_4357 = io_in_bits_DecodeIn_data_src2[56] ? io_in_bits_DecodeIn_data_src1[56] : io_in_bits_DecodeIn_data_src3[
    56]; // @[PALU.scala 477:46]
  wire  _T_4362 = io_in_bits_DecodeIn_data_src2[57] ? io_in_bits_DecodeIn_data_src1[57] : io_in_bits_DecodeIn_data_src3[
    57]; // @[PALU.scala 477:46]
  wire  _T_4367 = io_in_bits_DecodeIn_data_src2[58] ? io_in_bits_DecodeIn_data_src1[58] : io_in_bits_DecodeIn_data_src3[
    58]; // @[PALU.scala 477:46]
  wire  _T_4372 = io_in_bits_DecodeIn_data_src2[59] ? io_in_bits_DecodeIn_data_src1[59] : io_in_bits_DecodeIn_data_src3[
    59]; // @[PALU.scala 477:46]
  wire  _T_4377 = io_in_bits_DecodeIn_data_src2[60] ? io_in_bits_DecodeIn_data_src1[60] : io_in_bits_DecodeIn_data_src3[
    60]; // @[PALU.scala 477:46]
  wire  _T_4382 = io_in_bits_DecodeIn_data_src2[61] ? io_in_bits_DecodeIn_data_src1[61] : io_in_bits_DecodeIn_data_src3[
    61]; // @[PALU.scala 477:46]
  wire  _T_4387 = io_in_bits_DecodeIn_data_src2[62] ? io_in_bits_DecodeIn_data_src1[62] : io_in_bits_DecodeIn_data_src3[
    62]; // @[PALU.scala 477:46]
  wire  _T_4392 = io_in_bits_DecodeIn_data_src2[63] ? io_in_bits_DecodeIn_data_src1[63] : io_in_bits_DecodeIn_data_src3[
    63]; // @[PALU.scala 477:46]
  wire [9:0] _T_4401 = {_T_4077,_T_4082,_T_4087,_T_4092,_T_4097,_T_4102,_T_4107,_T_4112,_T_4117,_T_4122}; // @[Cat.scala 30:58]
  wire [18:0] _T_4410 = {_T_4401,_T_4127,_T_4132,_T_4137,_T_4142,_T_4147,_T_4152,_T_4157,_T_4162,_T_4167}; // @[Cat.scala 30:58]
  wire [27:0] _T_4419 = {_T_4410,_T_4172,_T_4177,_T_4182,_T_4187,_T_4192,_T_4197,_T_4202,_T_4207,_T_4212}; // @[Cat.scala 30:58]
  wire [36:0] _T_4428 = {_T_4419,_T_4217,_T_4222,_T_4227,_T_4232,_T_4237,_T_4242,_T_4247,_T_4252,_T_4257}; // @[Cat.scala 30:58]
  wire [45:0] _T_4437 = {_T_4428,_T_4262,_T_4267,_T_4272,_T_4277,_T_4282,_T_4287,_T_4292,_T_4297,_T_4302}; // @[Cat.scala 30:58]
  wire [54:0] _T_4446 = {_T_4437,_T_4307,_T_4312,_T_4317,_T_4322,_T_4327,_T_4332,_T_4337,_T_4342,_T_4347}; // @[Cat.scala 30:58]
  wire [63:0] _T_4455 = {_T_4446,_T_4352,_T_4357,_T_4362,_T_4367,_T_4372,_T_4377,_T_4382,_T_4387,_T_4392}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_825 = {{32'd0}, _T_4455[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4529 = _GEN_825 & 64'hffffffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4531 = {_T_4455[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4533 = _T_4531 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4534 = _T_4529 | _T_4533; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_826 = {{16'd0}, _T_4534[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4539 = _GEN_826 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4541 = {_T_4534[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4543 = _T_4541 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4544 = _T_4539 | _T_4543; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_827 = {{8'd0}, _T_4544[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4549 = _GEN_827 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4551 = {_T_4544[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4553 = _T_4551 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4554 = _T_4549 | _T_4553; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_828 = {{4'd0}, _T_4554[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4559 = _GEN_828 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4561 = {_T_4554[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4563 = _T_4561 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4564 = _T_4559 | _T_4563; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_829 = {{2'd0}, _T_4564[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4569 = _GEN_829 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4571 = {_T_4564[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4573 = _T_4571 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4574 = _T_4569 | _T_4573; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_830 = {{1'd0}, _T_4574[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4579 = _GEN_830 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4581 = {_T_4574[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4583 = _T_4581 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4584 = _T_4579 | _T_4583; // @[Bitwise.scala 103:39]
  wire [63:0] cmixRes = io_in_bits_Pctrl_isCmix ? _T_4584 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 598:17 599:17]
  wire [7:0] _GEN_610 = 3'h0 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[7:0]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_611 = 3'h1 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[15:8]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_612 = 3'h2 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[23:16]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_613 = 3'h3 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[31:24]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_614 = 3'h4 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[39:32]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_615 = 3'h5 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[47:40]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_616 = 3'h6 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[55:48]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_617 = 3'h7 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[63:56]; // @[PALU.scala 485:31 486:21]
  wire [63:0] _T_4679 = {_GEN_617,_GEN_616,_GEN_615,_GEN_614,_GEN_613,_GEN_612,_GEN_611,_GEN_610}; // @[Cat.scala 30:58]
  wire [63:0] insbRes = io_in_bits_Pctrl_isInsertb ? _T_4679 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 604:20 605:17]
  wire [31:0] _T_4683 = io_in_bits_Pctrl_isPackbb | io_in_bits_Pctrl_isPacktb ? io_in_bits_DecodeIn_data_src2[31:0] :
    io_in_bits_DecodeIn_data_src2[63:32]; // @[PALU.scala 611:25]
  wire [31:0] _T_4687 = io_in_bits_Pctrl_isPackbb | io_in_bits_Pctrl_isPackbt ? io_in_bits_DecodeIn_data_src1[31:0] :
    io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 612:25]
  wire [63:0] _T_4689 = {_T_4683,_T_4687}; // @[Cat.scala 30:58]
  wire [63:0] _T_4690 = {_T_4687,_T_4683}; // @[Cat.scala 30:58]
  wire [63:0] _T_4691 = io_in_bits_Pctrl_isPackbb | io_in_bits_Pctrl_isPacktt ? _T_4689 : _T_4690; // @[PALU.scala 613:23]
  wire [63:0] packRes = io_in_bits_Pctrl_isPack ? _T_4691 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 610:17 613:17]
  wire [63:0] _GEN_620 = io_in_bits_Pctrl_isInsertb ? insbRes : adderRes_final; // @[PALU.scala 655:26 656:28 659:28]
  wire  _GEN_621 = io_in_bits_Pctrl_isInsertb ? 1'h0 : adderOV; // @[PALU.scala 655:26 657:39 660:39]
  wire [63:0] _GEN_622 = io_in_bits_Pctrl_isBitrev ? bitrevRes : _GEN_620; // @[PALU.scala 652:25 653:28]
  wire  _GEN_623 = io_in_bits_Pctrl_isBitrev ? 1'h0 : _GEN_621; // @[PALU.scala 652:25 654:39]
  wire [63:0] _GEN_624 = io_in_bits_Pctrl_isPbs ? pbsRes : _GEN_622; // @[PALU.scala 649:22 650:28]
  wire  _GEN_625 = io_in_bits_Pctrl_isPbs ? 1'h0 : _GEN_623; // @[PALU.scala 649:22 651:39]
  wire [63:0] _GEN_626 = io_in_bits_Pctrl_isUnpack ? unpackRes : _GEN_624; // @[PALU.scala 646:25 647:28]
  wire  _GEN_627 = io_in_bits_Pctrl_isUnpack ? 1'h0 : _GEN_625; // @[PALU.scala 646:25 648:39]
  wire [63:0] _GEN_628 = io_in_bits_Pctrl_isCnt ? cntRes : _GEN_626; // @[PALU.scala 643:22 644:28]
  wire  _GEN_629 = io_in_bits_Pctrl_isCnt ? 1'h0 : _GEN_627; // @[PALU.scala 643:22 645:39]
  wire [63:0] _GEN_630 = io_in_bits_Pctrl_isSat ? satRes : _GEN_628; // @[PALU.scala 640:22 641:28]
  wire  _GEN_631 = io_in_bits_Pctrl_isSat ? satOV : _GEN_629; // @[PALU.scala 640:22 642:39]
  wire [63:0] _GEN_632 = io_in_bits_Pctrl_isClip ? clipRes : _GEN_630; // @[PALU.scala 637:23 638:28]
  wire  _GEN_633 = io_in_bits_Pctrl_isClip ? clipOV : _GEN_631; // @[PALU.scala 637:23 639:39]
  wire [63:0] _GEN_634 = io_in_bits_Pctrl_isCompare ? compareRes : _GEN_632; // @[PALU.scala 634:26 635:28]
  wire  _GEN_635 = io_in_bits_Pctrl_isCompare ? 1'h0 : _GEN_633; // @[PALU.scala 634:26 636:39]
  wire [63:0] _GEN_636 = io_in_bits_Pctrl_isShifter ? shifterRes : _GEN_634; // @[PALU.scala 631:26 632:28]
  wire  _GEN_637 = io_in_bits_Pctrl_isShifter ? shifterOV : _GEN_635; // @[PALU.scala 631:26 633:39]
  wire [63:0] _GEN_638 = io_in_bits_Pctrl_isAdder ? adderRes_final : _GEN_636; // @[PALU.scala 628:24 629:28]
  wire  _GEN_639 = io_in_bits_Pctrl_isAdder ? adderOV : _GEN_637; // @[PALU.scala 628:24 630:39]
  wire [63:0] _GEN_640 = io_in_bits_Pctrl_isCmix ? cmixRes : _GEN_638; // @[PALU.scala 625:23 626:28]
  wire  _GEN_641 = io_in_bits_Pctrl_isCmix ? 1'h0 : _GEN_639; // @[PALU.scala 625:23 627:39]
  wire [63:0] _GEN_642 = io_in_bits_Pctrl_isSwap ? swapRes : _GEN_640; // @[PALU.scala 622:23 623:28]
  wire  _GEN_643 = io_in_bits_Pctrl_isSwap ? 1'h0 : _GEN_641; // @[PALU.scala 622:23 624:39]
  wire [63:0] _GEN_644 = io_in_bits_Pctrl_isMaxMin ? maxminRes : _GEN_642; // @[PALU.scala 619:25 620:28]
  wire  _GEN_645 = io_in_bits_Pctrl_isMaxMin ? 1'h0 : _GEN_643; // @[PALU.scala 619:25 621:39]
  assign io_in_ready = ~io_in_valid | _T_1; // @[PALU.scala 37:27]
  assign io_out_valid = io_in_valid; // @[PALU.scala 38:17]
  assign io_out_bits_result = io_in_bits_Pctrl_isPack ? packRes : _GEN_644; // @[PALU.scala 616:17 617:28]
  assign io_out_bits_DecodeOut_cf_pc = io_in_bits_DecodeIn_cf_pc; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_cf_runahead_checkpoint_id = io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_ctrl_rfWen = io_in_bits_DecodeIn_ctrl_rfWen; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_ctrl_rfDest = io_in_bits_DecodeIn_ctrl_rfDest; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_pext_OV = io_in_bits_Pctrl_isPack ? 1'h0 : _GEN_645; // @[PALU.scala 616:17 618:39]
  assign io_out_bits_DecodeOut_InstNo = io_in_bits_DecodeIn_InstNo; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_InstFlag = io_in_bits_DecodeIn_InstFlag; // @[PALU.scala 39:27]
endmodule
module PMDU(
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_DecodeIn_cf_pc,
  input  [63:0]  io_in_bits_DecodeIn_cf_runahead_checkpoint_id,
  input  [6:0]   io_in_bits_DecodeIn_ctrl_fuOpType,
  input          io_in_bits_DecodeIn_ctrl_rfWen,
  input  [4:0]   io_in_bits_DecodeIn_ctrl_rfDest,
  input  [63:0]  io_in_bits_DecodeIn_data_src1,
  input  [63:0]  io_in_bits_DecodeIn_data_src2,
  input  [63:0]  io_in_bits_DecodeIn_data_src3,
  input  [4:0]   io_in_bits_DecodeIn_InstNo,
  input          io_in_bits_DecodeIn_InstFlag,
  input          io_in_bits_Pctrl_isMul_16,
  input          io_in_bits_Pctrl_isMul_8,
  input          io_in_bits_Pctrl_isMSW_3232,
  input          io_in_bits_Pctrl_isMSW_3216,
  input          io_in_bits_Pctrl_isS1632,
  input          io_in_bits_Pctrl_isS1664,
  input          io_in_bits_Pctrl_is832,
  input          io_in_bits_Pctrl_is3264,
  input          io_in_bits_Pctrl_is1664,
  input          io_in_bits_Pctrl_isQ15orQ31,
  input          io_in_bits_Pctrl_isC31,
  input          io_in_bits_Pctrl_isQ15_64ONLY,
  input          io_in_bits_Pctrl_isQ63_64ONLY,
  input          io_in_bits_Pctrl_isMul_32_64ONLY,
  input          io_in_bits_Pctrl_isPMA_64ONLY,
  input  [17:0]  io_in_bits_Pctrl_mulres9_0,
  input  [17:0]  io_in_bits_Pctrl_mulres9_1,
  input  [17:0]  io_in_bits_Pctrl_mulres9_2,
  input  [17:0]  io_in_bits_Pctrl_mulres9_3,
  input  [33:0]  io_in_bits_Pctrl_mulres17_0,
  input  [33:0]  io_in_bits_Pctrl_mulres17_1,
  input  [65:0]  io_in_bits_Pctrl_mulres33_0,
  input  [129:0] io_in_bits_Pctrl_mulres65_0,
  input          io_out_ready,
  output         io_out_valid,
  output [63:0]  io_out_bits_result,
  output [38:0]  io_out_bits_DecodeOut_cf_pc,
  output [63:0]  io_out_bits_DecodeOut_cf_runahead_checkpoint_id,
  output [6:0]   io_out_bits_DecodeOut_ctrl_fuOpType,
  output         io_out_bits_DecodeOut_ctrl_rfWen,
  output [4:0]   io_out_bits_DecodeOut_ctrl_rfDest,
  output [63:0]  io_out_bits_DecodeOut_data_src1,
  output [63:0]  io_out_bits_DecodeOut_data_src2,
  output [63:0]  io_out_bits_DecodeOut_data_src3,
  output         io_out_bits_DecodeOut_pext_OV,
  output [4:0]   io_out_bits_DecodeOut_InstNo,
  output         io_out_bits_DecodeOut_InstFlag,
  output         io_FirstStageFire
);
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [32:0] _T_718 = {io_out_bits_DecodeOut_data_src3[63],io_out_bits_DecodeOut_data_src3[63:32]}; // @[Cat.scala 30:58]
  wire [1:0] _T_1035 = io_out_bits_DecodeOut_data_src3[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1036 = {_T_1035,io_out_bits_DecodeOut_data_src3[63:32]}; // @[Cat.scala 30:58]
  wire  _T_467 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h4; // @[PMDU.scala 849:59]
  wire [31:0] _T_469 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h4 ? io_out_bits_DecodeOut_data_src3[63:32] : 32'h0
    ; // @[PMDU.scala 849:45]
  wire [32:0] _T_471 = {_T_469[31],_T_469}; // @[Cat.scala 30:58]
  wire [33:0] _GEN_88 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _T_471} : 34'h0; // @[PMDU.scala 836:50 865:34]
  wire [33:0] _GEN_101 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_88; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_113 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_101; // @[PMDU.scala 735:40]
  wire [33:0] _GEN_223 = io_in_bits_Pctrl_is832 ? {{2'd0}, io_out_bits_DecodeOut_data_src3[63:32]} : _GEN_113; // @[PMDU.scala 1051:39 1078:30]
  wire [33:0] _GEN_244 = io_in_bits_Pctrl_isS1664 ? _GEN_113 : _GEN_223; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_257 = io_in_bits_Pctrl_isS1632 ? _T_1036 : _GEN_244; // @[PMDU.scala 1000:41 1020:30]
  wire [33:0] _GEN_273 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_718} : _GEN_257; // @[PMDU.scala 963:44 979:30]
  wire [33:0] adder34_0_1 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_718} : _GEN_273; // @[PMDU.scala 929:38 938:30]
  wire [32:0] _T_638 = {io_out_bits_DecodeOut_data_src3[31],io_out_bits_DecodeOut_data_src3[31:0]}; // @[Cat.scala 30:58]
  wire [1:0] _T_968 = io_out_bits_DecodeOut_data_src3[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_969 = {_T_968,io_out_bits_DecodeOut_data_src3[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_417 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h4 ? io_out_bits_DecodeOut_data_src3[31:0] : 32'h0; // @[PMDU.scala 849:45]
  wire [32:0] _T_419 = {_T_417[31],_T_417}; // @[Cat.scala 30:58]
  wire [33:0] _GEN_85 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _T_419} : 34'h0; // @[PMDU.scala 836:50 865:34]
  wire [33:0] _GEN_98 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_85; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_110 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_98; // @[PMDU.scala 735:40]
  wire [33:0] _GEN_218 = io_in_bits_Pctrl_is832 ? {{2'd0}, io_out_bits_DecodeOut_data_src3[31:0]} : _GEN_110; // @[PMDU.scala 1051:39 1078:30]
  wire [33:0] _GEN_239 = io_in_bits_Pctrl_isS1664 ? _GEN_110 : _GEN_218; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_252 = io_in_bits_Pctrl_isS1632 ? _T_969 : _GEN_239; // @[PMDU.scala 1000:41 1020:30]
  wire [33:0] _GEN_270 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_638} : _GEN_252; // @[PMDU.scala 963:44 979:30]
  wire [33:0] adder34_0_0 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_638} : _GEN_270; // @[PMDU.scala 929:38 938:30]
  wire [70:0] _T_12 = {adder34_0_1,3'h0,adder34_0_0}; // @[Cat.scala 30:58]
  wire [64:0] _T_512 = {io_out_bits_DecodeOut_data_src3[63],io_out_bits_DecodeOut_data_src3}; // @[Cat.scala 30:58]
  wire  _T_533 = ~(_T_467 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h1d); // @[PMDU.scala 904:31]
  wire [1:0] _T_555 = io_out_bits_DecodeOut_data_src3[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_556 = {_T_555,io_out_bits_DecodeOut_data_src3}; // @[Cat.scala 30:58]
  wire [65:0] _T_557 = _T_533 ? _T_556 : 66'h0; // @[PMDU.scala 908:33]
  wire [70:0] _GEN_66 = io_in_bits_Pctrl_isPMA_64ONLY ? {{5'd0}, _T_557} : _T_12; // @[PMDU.scala 728:15 902:50 908:27]
  wire [70:0] _GEN_72 = io_in_bits_Pctrl_isQ63_64ONLY ? {{6'd0}, _T_512} : _GEN_66; // @[PMDU.scala 886:50 888:27]
  wire [70:0] _GEN_79 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_12 : _GEN_72; // @[PMDU.scala 728:15 884:53]
  wire [70:0] _GEN_92 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_12 : _GEN_79; // @[PMDU.scala 728:15 836:50]
  wire [70:0] _GEN_104 = io_in_bits_Pctrl_isMul_8 ? _T_12 : _GEN_92; // @[PMDU.scala 728:15 779:45]
  wire [70:0] _GEN_116 = io_in_bits_Pctrl_isMul_16 ? _T_12 : _GEN_104; // @[PMDU.scala 728:15 735:40]
  wire  _T_1198 = ~io_out_bits_DecodeOut_ctrl_fuOpType[4]; // @[PMDU.scala 1090:24]
  wire [65:0] _T_1216 = {2'h0,io_out_bits_DecodeOut_data_src3}; // @[Cat.scala 30:58]
  wire [65:0] _GEN_176 = _T_1198 ? _T_556 : _T_1216; // @[PMDU.scala 676:24 677:15 679:15]
  wire [31:0] _T_1413 = io_out_bits_DecodeOut_ctrl_fuOpType[4] ? 32'h0 : io_out_bits_DecodeOut_data_src3[31:0]; // @[PMDU.scala 1186:29]
  wire [70:0] _GEN_195 = io_in_bits_Pctrl_isC31 ? {{39'd0}, _T_1413} : _GEN_116; // @[PMDU.scala 1183:39 1186:23]
  wire [70:0] _GEN_200 = io_in_bits_Pctrl_isQ15orQ31 ? {{38'd0}, _T_638} : _GEN_195; // @[PMDU.scala 1149:44 1167:23]
  wire [70:0] _GEN_204 = io_in_bits_Pctrl_is1664 ? {{7'd0}, io_out_bits_DecodeOut_data_src3} : _GEN_200; // @[PMDU.scala 1126:40 1136:23]
  wire [70:0] _GEN_211 = io_in_bits_Pctrl_is3264 ? {{5'd0}, _GEN_176} : _GEN_204; // @[PMDU.scala 1089:40 1098:23]
  wire [70:0] _GEN_229 = io_in_bits_Pctrl_is832 ? _GEN_116 : _GEN_211; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_235 = io_in_bits_Pctrl_isS1664 ? {{7'd0}, io_out_bits_DecodeOut_data_src1} : _GEN_229; // @[PMDU.scala 1046:41 1047:19]
  wire [70:0] _GEN_262 = io_in_bits_Pctrl_isS1632 ? _GEN_116 : _GEN_235; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_279 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_116 : _GEN_262; // @[PMDU.scala 963:44]
  wire [70:0] adder68_0 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_116 : _GEN_279; // @[PMDU.scala 929:38]
  wire  _T_686 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h1; // @[PMDU.scala 933:69]
  wire  _T_687 = io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h2 & io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h1; // @[PMDU.scala 933:52]
  wire [32:0] _T_720 = _T_687 ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire  _T_694 = io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h3; // @[PMDU.scala 935:40]
  wire  _T_697 = io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h3 & _T_686; // @[PMDU.scala 935:52]
  wire [32:0] _T_703 = io_in_bits_Pctrl_mulres65_0[63:31] + 33'h1; // @[PMDU.scala 936:164]
  wire [32:0] _T_705 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_703 : io_in_bits_Pctrl_mulres65_0[63:31]; // @[PMDU.scala 936:41]
  wire [33:0] _T_711 = io_in_bits_Pctrl_mulres65_0[63:30] + 34'h1; // @[PMDU.scala 937:164]
  wire [33:0] _T_713 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_711 : io_in_bits_Pctrl_mulres65_0[63:30]; // @[PMDU.scala 937:41]
  wire [31:0] _T_715 = ~_T_697 ? _T_705[32:1] : _T_713[32:1]; // @[PMDU.scala 936:32]
  wire [32:0] _T_722 = {_T_715[31],_T_715}; // @[Cat.scala 30:58]
  wire [32:0] _T_723 = _T_720 ^ _T_722; // @[PMDU.scala 939:53]
  wire  _T_847 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h7; // @[PMDU.scala 968:41]
  wire  _T_880 = io_out_bits_DecodeOut_data_src1[63:32] == 32'h80000000; // @[PMDU.scala 975:62]
  wire  _T_855 = _T_694 | io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h5 | io_out_bits_DecodeOut_ctrl_fuOpType[6:4]
     == 3'h7; // @[PMDU.scala 969:93]
  wire [15:0] _T_858 = _T_855 ? io_out_bits_DecodeOut_data_src2[63:48] : io_out_bits_DecodeOut_data_src2[47:32]; // @[PMDU.scala 970:36]
  wire [32:0] _T_864 = io_in_bits_Pctrl_mulres65_0[47:15] + 33'h1; // @[PMDU.scala 971:165]
  wire [32:0] _T_866 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_864 : io_in_bits_Pctrl_mulres65_0[47:15]; // @[PMDU.scala 971:42]
  wire [32:0] _T_872 = io_in_bits_Pctrl_mulres65_0[46:14] + 33'h1; // @[PMDU.scala 972:164]
  wire [32:0] _T_874 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_872 : io_in_bits_Pctrl_mulres65_0[46:14]; // @[PMDU.scala 972:41]
  wire [31:0] _T_876 = ~_T_847 ? _T_866[32:1] : _T_874[32:1]; // @[PMDU.scala 971:33]
  wire [31:0] _GEN_146 = _T_847 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80000000 & _T_858 == 16'h8000 ? 32'h7fffffff
     : _T_876; // @[PMDU.scala 975:127 974:23 977:27]
  wire [32:0] _T_892 = {_GEN_146[31],_GEN_146}; // @[Cat.scala 30:58]
  wire  _T_934 = io_out_bits_DecodeOut_ctrl_fuOpType[6:1] == 6'h13; // @[PMDU.scala 1002:95]
  wire  _T_935 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h34 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h36 |
    io_out_bits_DecodeOut_ctrl_fuOpType[6:1] == 6'h13; // @[PMDU.scala 1002:78]
  wire [33:0] _T_1038 = _T_935 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_1041 = io_in_bits_Pctrl_mulres65_0[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1042 = {_T_1041,io_in_bits_Pctrl_mulres65_0[31:0]}; // @[Cat.scala 30:58]
  wire [33:0] _T_1043 = _T_1038 ^ _T_1042; // @[PMDU.scala 1021:57]
  wire  _T_402 = io_out_bits_DecodeOut_ctrl_fuOpType[4:3] == 2'h1; // @[PMDU.scala 838:40]
  wire  _T_404 = io_out_bits_DecodeOut_ctrl_fuOpType[4:3] == 2'h2; // @[PMDU.scala 839:40]
  wire [15:0] _T_460 = _T_404 ? io_out_bits_DecodeOut_data_src1[47:32] : io_out_bits_DecodeOut_data_src1[63:48]; // @[PMDU.scala 842:70]
  wire [15:0] _T_461 = _T_402 ? io_out_bits_DecodeOut_data_src1[47:32] : _T_460; // @[PMDU.scala 842:40]
  wire [15:0] _T_464 = _T_402 ? io_out_bits_DecodeOut_data_src2[47:32] : io_out_bits_DecodeOut_data_src2[63:48]; // @[PMDU.scala 843:40]
  wire  _T_476 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h6; // @[PMDU.scala 853:44]
  wire [30:0] _GEN_49 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h6 ? 31'h7fff : 31'h7fffffff; // @[PMDU.scala 853:57 854:36 856:36]
  wire [16:0] _T_482 = io_in_bits_Pctrl_mulres65_0[30] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_483 = {_T_482,io_in_bits_Pctrl_mulres65_0[30:15]}; // @[Cat.scala 30:58]
  wire [32:0] _T_485 = {io_in_bits_Pctrl_mulres65_0[31],io_in_bits_Pctrl_mulres65_0[31:0]}; // @[Cat.scala 30:58]
  wire [33:0] _T_486 = {_T_485, 1'h0}; // @[PMDU.scala 862:64]
  wire [32:0] _T_489 = {_T_486[31],_T_486[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_50 = _T_476 ? _T_483 : _T_489; // @[PMDU.scala 859:57 860:36 862:36]
  wire [32:0] _GEN_52 = _T_461 == 16'h8000 & _T_464 == 16'h8000 ? {{2'd0}, _GEN_49} : _GEN_50; // @[PMDU.scala 851:77]
  wire [33:0] _GEN_89 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _GEN_52} : 34'h0; // @[PMDU.scala 836:50 866:34]
  wire [33:0] _GEN_102 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_89; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_114 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_102; // @[PMDU.scala 735:40]
  wire  _T_1156 = ~_T_476; // @[PMDU.scala 1073:38]
  wire [14:0] _T_1160 = io_in_bits_Pctrl_mulres17_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1161 = {_T_1160,io_in_bits_Pctrl_mulres17_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1162 = {15'h0,io_in_bits_Pctrl_mulres17_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_170 = _T_1156 ? _T_1161 : _T_1162; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_224 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_170} : _GEN_114; // @[PMDU.scala 1051:39 1079:30]
  wire [33:0] _GEN_245 = io_in_bits_Pctrl_isS1664 ? _GEN_114 : _GEN_224; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_258 = io_in_bits_Pctrl_isS1632 ? _T_1043 : _GEN_245; // @[PMDU.scala 1000:41 1021:30]
  wire [33:0] _GEN_274 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_892} : _GEN_258; // @[PMDU.scala 963:44 980:30]
  wire [33:0] adder34_1_1 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_723} : _GEN_274; // @[PMDU.scala 929:38 939:30]
  wire [32:0] _T_623 = io_in_bits_Pctrl_mulres33_0[63:31] + 33'h1; // @[PMDU.scala 936:120]
  wire [32:0] _T_625 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_623 : io_in_bits_Pctrl_mulres33_0[63:31]; // @[PMDU.scala 936:41]
  wire [33:0] _T_631 = io_in_bits_Pctrl_mulres33_0[63:30] + 34'h1; // @[PMDU.scala 937:120]
  wire [33:0] _T_633 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_631 : io_in_bits_Pctrl_mulres33_0[63:30]; // @[PMDU.scala 937:41]
  wire [31:0] _T_635 = ~_T_697 ? _T_625[32:1] : _T_633[32:1]; // @[PMDU.scala 936:32]
  wire [32:0] _T_642 = {_T_635[31],_T_635}; // @[Cat.scala 30:58]
  wire [32:0] _T_643 = _T_720 ^ _T_642; // @[PMDU.scala 939:53]
  wire  _T_803 = io_out_bits_DecodeOut_data_src1[31:0] == 32'h80000000; // @[PMDU.scala 975:62]
  wire [15:0] _T_781 = _T_855 ? io_out_bits_DecodeOut_data_src2[31:16] : io_out_bits_DecodeOut_data_src2[15:0]; // @[PMDU.scala 970:36]
  wire [32:0] _T_787 = io_in_bits_Pctrl_mulres33_0[47:15] + 33'h1; // @[PMDU.scala 971:121]
  wire [32:0] _T_789 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_787 : io_in_bits_Pctrl_mulres33_0[47:15]; // @[PMDU.scala 971:42]
  wire [32:0] _T_795 = io_in_bits_Pctrl_mulres33_0[46:14] + 33'h1; // @[PMDU.scala 972:120]
  wire [32:0] _T_797 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_795 : io_in_bits_Pctrl_mulres33_0[46:14]; // @[PMDU.scala 972:41]
  wire [31:0] _T_799 = ~_T_847 ? _T_789[32:1] : _T_797[32:1]; // @[PMDU.scala 971:33]
  wire [31:0] _GEN_139 = _T_847 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80000000 & _T_781 == 16'h8000 ? 32'h7fffffff
     : _T_799; // @[PMDU.scala 975:127 974:23 977:27]
  wire [32:0] _T_815 = {_GEN_139[31],_GEN_139}; // @[Cat.scala 30:58]
  wire  _T_922 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h5; // @[PMDU.scala 1001:61]
  wire  _T_924 = io_out_bits_DecodeOut_ctrl_fuOpType[6:5] == 2'h1; // @[PMDU.scala 1001:91]
  wire  _T_929 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] < 4'h3 | io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h5 &
    io_out_bits_DecodeOut_ctrl_fuOpType[6:5] == 2'h1 & io_out_bits_DecodeOut_ctrl_fuOpType[4:3] != 2'h0; // @[PMDU.scala 1001:44]
  wire [31:0] _T_962 = _T_929 ? io_in_bits_Pctrl_mulres33_0[31:0] : io_in_bits_Pctrl_mulres17_1[31:0]; // @[PMDU.scala 1011:39]
  wire [1:0] _T_974 = _T_962[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_975 = {_T_974,_T_962}; // @[Cat.scala 30:58]
  wire [33:0] _T_976 = _T_1038 ^ _T_975; // @[PMDU.scala 1021:57]
  wire [15:0] _T_408 = _T_404 ? io_out_bits_DecodeOut_data_src1[15:0] : io_out_bits_DecodeOut_data_src1[31:16]; // @[PMDU.scala 842:70]
  wire [15:0] _T_409 = _T_402 ? io_out_bits_DecodeOut_data_src1[15:0] : _T_408; // @[PMDU.scala 842:40]
  wire [15:0] _T_412 = _T_402 ? io_out_bits_DecodeOut_data_src2[15:0] : io_out_bits_DecodeOut_data_src2[31:16]; // @[PMDU.scala 843:40]
  wire  _T_422 = _T_409 == 16'h8000 & _T_412 == 16'h8000; // @[PMDU.scala 851:50]
  wire [16:0] _T_430 = io_in_bits_Pctrl_mulres33_0[30] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_431 = {_T_430,io_in_bits_Pctrl_mulres33_0[30:15]}; // @[Cat.scala 30:58]
  wire [32:0] _T_433 = {io_in_bits_Pctrl_mulres33_0[31],io_in_bits_Pctrl_mulres33_0[31:0]}; // @[Cat.scala 30:58]
  wire [33:0] _T_434 = {_T_433, 1'h0}; // @[PMDU.scala 862:64]
  wire [32:0] _T_437 = {_T_434[31],_T_434[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_41 = _T_476 ? _T_431 : _T_437; // @[PMDU.scala 859:57 860:36 862:36]
  wire [32:0] _GEN_43 = _T_409 == 16'h8000 & _T_412 == 16'h8000 ? {{2'd0}, _GEN_49} : _GEN_41; // @[PMDU.scala 851:77]
  wire [33:0] _GEN_86 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _GEN_43} : 34'h0; // @[PMDU.scala 836:50 866:34]
  wire [33:0] _GEN_99 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_86; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_111 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_99; // @[PMDU.scala 735:40]
  wire [14:0] _T_1121 = io_in_bits_Pctrl_mulres9_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1122 = {_T_1121,io_in_bits_Pctrl_mulres9_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1123 = {15'h0,io_in_bits_Pctrl_mulres9_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_166 = _T_1156 ? _T_1122 : _T_1123; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_219 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_166} : _GEN_111; // @[PMDU.scala 1051:39 1079:30]
  wire [33:0] _GEN_240 = io_in_bits_Pctrl_isS1664 ? _GEN_111 : _GEN_219; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_253 = io_in_bits_Pctrl_isS1632 ? _T_976 : _GEN_240; // @[PMDU.scala 1000:41 1021:30]
  wire [33:0] _GEN_271 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_815} : _GEN_253; // @[PMDU.scala 963:44 980:30]
  wire [33:0] adder34_1_0 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_643} : _GEN_271; // @[PMDU.scala 929:38 939:30]
  wire [70:0] _T_13 = {adder34_1_1,3'h0,adder34_1_0}; // @[Cat.scala 30:58]
  wire [64:0] _T_515 = {io_in_bits_Pctrl_mulres65_0[63],io_in_bits_Pctrl_mulres65_0[63:0]}; // @[Cat.scala 30:58]
  wire  _T_538 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h5 | io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h7; // @[PMDU.scala 905:59]
  wire  _T_541 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h5 | io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h7 |
    _T_934; // @[PMDU.scala 905:90]
  wire [65:0] _T_559 = _T_541 ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_563 = io_in_bits_Pctrl_mulres33_0[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_564 = {_T_563,io_in_bits_Pctrl_mulres33_0[63:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_565 = _T_559 ^ _T_564; // @[PMDU.scala 909:47]
  wire [70:0] _GEN_67 = io_in_bits_Pctrl_isPMA_64ONLY ? {{5'd0}, _T_565} : _T_13; // @[PMDU.scala 729:15 902:50 909:27]
  wire [70:0] _GEN_73 = io_in_bits_Pctrl_isQ63_64ONLY ? {{6'd0}, _T_515} : _GEN_67; // @[PMDU.scala 886:50 889:27]
  wire [70:0] _GEN_80 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_13 : _GEN_73; // @[PMDU.scala 729:15 884:53]
  wire [70:0] _GEN_93 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_13 : _GEN_80; // @[PMDU.scala 729:15 836:50]
  wire [70:0] _GEN_105 = io_in_bits_Pctrl_isMul_8 ? _T_13 : _GEN_93; // @[PMDU.scala 729:15 779:45]
  wire [70:0] _GEN_117 = io_in_bits_Pctrl_isMul_16 ? _T_13 : _GEN_105; // @[PMDU.scala 729:15 735:40]
  wire [31:0] _T_1107 = io_in_bits_Pctrl_mulres65_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1108 = {_T_1107,io_in_bits_Pctrl_mulres65_0[31:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1218 = io_out_bits_DecodeOut_ctrl_fuOpType[0] ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_1205 = {io_in_bits_Pctrl_mulres33_0[64],io_in_bits_Pctrl_mulres33_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1206 = {1'h0,io_in_bits_Pctrl_mulres33_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _GEN_174 = _T_1198 ? _T_1205 : _T_1206; // @[PMDU.scala 676:24 677:15 679:15]
  wire [65:0] _T_1219 = _T_1218 ^ _GEN_174; // @[PMDU.scala 1099:41]
  wire  _T_1258 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h56; // @[PMDU.scala 1128:90]
  wire  _T_1260 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h5e; // @[PMDU.scala 1128:119]
  wire  _T_1261 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h45 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h55 |
    io_out_bits_DecodeOut_ctrl_fuOpType == 7'h56 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h5e; // @[PMDU.scala 1128:107]
  wire [63:0] _T_1279 = _T_1261 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1269 = _T_467 ? io_in_bits_Pctrl_mulres33_0[31:0] : io_in_bits_Pctrl_mulres17_0[31:0]; // @[PMDU.scala 1132:23]
  wire [31:0] _T_1282 = _T_1269[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1283 = {_T_1282,_T_1269}; // @[Cat.scala 30:58]
  wire [63:0] _T_1284 = _T_1279 ^ _T_1283; // @[PMDU.scala 1137:50]
  wire [1:0] _T_1285 = {_T_1261,1'h0}; // @[Cat.scala 30:58]
  wire  _T_1266 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h4d | _T_1258 | _T_1260; // @[PMDU.scala 1129:78]
  wire [1:0] _T_1286 = {_T_1266,1'h0}; // @[Cat.scala 30:58]
  wire [2:0] _T_1287 = _T_1285 + _T_1286; // @[PMDU.scala 1137:101]
  wire [63:0] _GEN_303 = {{61'd0}, _T_1287}; // @[PMDU.scala 1137:69]
  wire [63:0] _T_1289 = _T_1284 + _GEN_303; // @[PMDU.scala 1137:69]
  wire  _T_1344 = _T_686 ? _T_402 : io_out_bits_DecodeOut_ctrl_fuOpType[4:3] == 2'h0; // @[PMDU.scala 1154:25]
  wire  _T_1349 = _T_686 ? _T_404 : _T_402; // @[PMDU.scala 1155:25]
  wire [15:0] _T_1353 = _T_1349 ? io_out_bits_DecodeOut_data_src1[15:0] : io_out_bits_DecodeOut_data_src1[31:16]; // @[PMDU.scala 1156:55]
  wire [15:0] _T_1354 = _T_1344 ? io_out_bits_DecodeOut_data_src1[15:0] : _T_1353; // @[PMDU.scala 1156:33]
  wire [15:0] _T_1357 = _T_1344 ? io_out_bits_DecodeOut_data_src2[15:0] : io_out_bits_DecodeOut_data_src2[31:16]; // @[PMDU.scala 1157:33]
  wire [63:0] _T_1364 = _T_476 ? 64'h7fff : 64'h7fffffff; // @[PMDU.scala 1163:28]
  wire [31:0] _T_1365 = io_in_bits_Pctrl_mulres65_0[31:0]; // @[PMDU.scala 1165:48]
  wire [16:0] _T_1367 = _T_1365[31:15]; // @[PMDU.scala 1165:62]
  wire [46:0] _T_1370 = _T_1367[16] ? 47'h7fffffffffff : 47'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1371 = {_T_1370,_T_1367}; // @[Cat.scala 30:58]
  wire [32:0] _T_1372 = {io_in_bits_Pctrl_mulres65_0[31:0], 1'h0}; // @[PMDU.scala 1165:87]
  wire [30:0] _T_1375 = _T_1372[32] ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1376 = {_T_1375,_T_1372}; // @[Cat.scala 30:58]
  wire [63:0] _T_1377 = _T_476 ? _T_1371 : _T_1376; // @[PMDU.scala 1165:28]
  wire [63:0] _GEN_189 = _T_1354 == 16'h8000 & _T_1357 == 16'h8000 ? _T_1364 : _T_1377; // @[PMDU.scala 1161:70 1163:22 1165:22]
  wire [32:0] _T_1383 = {_GEN_189[31],_GEN_189[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1418 = io_out_bits_DecodeOut_ctrl_fuOpType[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1420 = _T_1418 ^ io_in_bits_Pctrl_mulres65_0[31:0]; // @[PMDU.scala 1187:74]
  wire [63:0] _T_1421 = io_out_bits_DecodeOut_ctrl_fuOpType[4] ? io_in_bits_Pctrl_mulres65_0[63:0] : {{32'd0}, _T_1420}; // @[PMDU.scala 1187:29]
  wire [70:0] _GEN_196 = io_in_bits_Pctrl_isC31 ? {{7'd0}, _T_1421} : _GEN_117; // @[PMDU.scala 1183:39 1187:23]
  wire [70:0] _GEN_201 = io_in_bits_Pctrl_isQ15orQ31 ? {{38'd0}, _T_1383} : _GEN_196; // @[PMDU.scala 1149:44 1168:23]
  wire [70:0] _GEN_205 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1289} : _GEN_201; // @[PMDU.scala 1126:40 1137:23]
  wire [70:0] _GEN_212 = io_in_bits_Pctrl_is3264 ? {{5'd0}, _T_1219} : _GEN_205; // @[PMDU.scala 1089:40 1099:23]
  wire [70:0] _GEN_230 = io_in_bits_Pctrl_is832 ? _GEN_117 : _GEN_212; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_236 = io_in_bits_Pctrl_isS1664 ? {{7'd0}, _T_1108} : _GEN_230; // @[PMDU.scala 1046:41 1048:19]
  wire [70:0] _GEN_263 = io_in_bits_Pctrl_isS1632 ? _GEN_117 : _GEN_236; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_280 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_117 : _GEN_263; // @[PMDU.scala 963:44]
  wire [70:0] adder68_1 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_117 : _GEN_280; // @[PMDU.scala 929:38]
  wire [70:0] _T_5 = adder68_0 + adder68_1; // @[PMDU.scala 726:24]
  wire  _T_949 = _T_538 & (_T_467 | _T_476) | _T_934; // @[PMDU.scala 1003:146]
  wire [33:0] _T_1045 = _T_949 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1031 = _T_929 ? 32'h0 : io_in_bits_Pctrl_mulres33_0[31:0]; // @[PMDU.scala 1016:102]
  wire [1:0] _T_1048 = _T_1031[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1049 = {_T_1048,_T_1031}; // @[Cat.scala 30:58]
  wire [33:0] _T_1050 = _T_1045 ^ _T_1049; // @[PMDU.scala 1022:56]
  wire [14:0] _T_1167 = io_in_bits_Pctrl_mulres17_1[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1168 = {_T_1167,io_in_bits_Pctrl_mulres17_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1169 = {15'h0,io_in_bits_Pctrl_mulres17_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_171 = _T_1156 ? _T_1168 : _T_1169; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_225 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_171} : 34'h0; // @[PMDU.scala 1051:39 1080:30]
  wire [33:0] _GEN_246 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_225; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_259 = io_in_bits_Pctrl_isS1632 ? _T_1050 : _GEN_246; // @[PMDU.scala 1000:41 1022:30]
  wire [33:0] _GEN_275 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_259; // @[PMDU.scala 963:44 981:30]
  wire [33:0] adder34_2_1 = io_in_bits_Pctrl_isMSW_3232 ? {{33'd0}, _T_687} : _GEN_275; // @[PMDU.scala 929:38 940:30]
  wire [31:0] _T_964 = _T_929 ? 32'h0 : io_in_bits_Pctrl_mulres17_0[31:0]; // @[PMDU.scala 1016:39]
  wire [1:0] _T_981 = _T_964[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_982 = {_T_981,_T_964}; // @[Cat.scala 30:58]
  wire [33:0] _T_983 = _T_1045 ^ _T_982; // @[PMDU.scala 1022:56]
  wire [14:0] _T_1128 = io_in_bits_Pctrl_mulres9_1[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1129 = {_T_1128,io_in_bits_Pctrl_mulres9_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1130 = {15'h0,io_in_bits_Pctrl_mulres9_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_167 = _T_1156 ? _T_1129 : _T_1130; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_220 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_167} : 34'h0; // @[PMDU.scala 1051:39 1080:30]
  wire [33:0] _GEN_241 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_220; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_254 = io_in_bits_Pctrl_isS1632 ? _T_983 : _GEN_241; // @[PMDU.scala 1000:41 1022:30]
  wire [33:0] _GEN_272 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_254; // @[PMDU.scala 963:44 981:30]
  wire [33:0] adder34_2_0 = io_in_bits_Pctrl_isMSW_3232 ? {{33'd0}, _T_687} : _GEN_272; // @[PMDU.scala 929:38 940:30]
  wire [70:0] _T_14 = {adder34_2_1,3'h0,adder34_2_0}; // @[Cat.scala 30:58]
  wire  _T_546 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h6 | _T_934; // @[PMDU.scala 906:59]
  wire [65:0] _T_567 = _T_546 ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_571 = io_in_bits_Pctrl_mulres65_0[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_572 = {_T_571,io_in_bits_Pctrl_mulres65_0[63:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_573 = _T_567 ^ _T_572; // @[PMDU.scala 910:47]
  wire [70:0] _GEN_68 = io_in_bits_Pctrl_isPMA_64ONLY ? {{5'd0}, _T_573} : _T_14; // @[PMDU.scala 730:15 902:50 910:27]
  wire [70:0] _GEN_74 = io_in_bits_Pctrl_isQ63_64ONLY ? 71'h0 : _GEN_68; // @[PMDU.scala 886:50 890:27]
  wire [70:0] _GEN_81 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_14 : _GEN_74; // @[PMDU.scala 730:15 884:53]
  wire [70:0] _GEN_94 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_14 : _GEN_81; // @[PMDU.scala 730:15 836:50]
  wire [70:0] _GEN_106 = io_in_bits_Pctrl_isMul_8 ? _T_14 : _GEN_94; // @[PMDU.scala 730:15 779:45]
  wire [70:0] _GEN_118 = io_in_bits_Pctrl_isMul_16 ? _T_14 : _GEN_106; // @[PMDU.scala 730:15 735:40]
  wire [31:0] _T_1112 = io_in_bits_Pctrl_mulres33_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1113 = {_T_1112,io_in_bits_Pctrl_mulres33_0[31:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1209 = {io_in_bits_Pctrl_mulres65_0[64],io_in_bits_Pctrl_mulres65_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1210 = {1'h0,io_in_bits_Pctrl_mulres65_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _GEN_175 = _T_1198 ? _T_1209 : _T_1210; // @[PMDU.scala 676:24 677:15 679:15]
  wire [65:0] _T_1222 = _T_1218 ^ _GEN_175; // @[PMDU.scala 1100:41]
  wire [31:0] _T_1274 = _T_467 ? 32'h0 : io_in_bits_Pctrl_mulres33_0[31:0]; // @[PMDU.scala 1134:23]
  wire [31:0] _T_1294 = _T_1274[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1295 = {_T_1294,_T_1274}; // @[Cat.scala 30:58]
  wire [63:0] _T_1296 = _T_1279 ^ _T_1295; // @[PMDU.scala 1138:50]
  wire [70:0] _GEN_197 = io_in_bits_Pctrl_isC31 ? {{70'd0}, io_out_bits_DecodeOut_ctrl_fuOpType[0]} : _GEN_118; // @[PMDU.scala 1183:39 1188:23]
  wire [70:0] _GEN_203 = io_in_bits_Pctrl_isQ15orQ31 ? _GEN_118 : _GEN_197; // @[PMDU.scala 1149:44]
  wire [70:0] _GEN_206 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1296} : _GEN_203; // @[PMDU.scala 1126:40 1138:23]
  wire [70:0] _GEN_213 = io_in_bits_Pctrl_is3264 ? {{5'd0}, _T_1222} : _GEN_206; // @[PMDU.scala 1089:40 1100:23]
  wire [70:0] _GEN_231 = io_in_bits_Pctrl_is832 ? _GEN_118 : _GEN_213; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_237 = io_in_bits_Pctrl_isS1664 ? {{7'd0}, _T_1113} : _GEN_231; // @[PMDU.scala 1046:41 1049:19]
  wire [70:0] _GEN_264 = io_in_bits_Pctrl_isS1632 ? _GEN_118 : _GEN_237; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_281 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_118 : _GEN_264; // @[PMDU.scala 963:44]
  wire [70:0] adder68_2 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_118 : _GEN_281; // @[PMDU.scala 929:38]
  wire [70:0] _T_7 = _T_5 + adder68_2; // @[PMDU.scala 726:36]
  wire [1:0] _T_1051 = _T_935 + _T_949; // @[PMDU.scala 1023:49]
  wire [14:0] _T_1174 = io_in_bits_Pctrl_mulres33_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1175 = {_T_1174,io_in_bits_Pctrl_mulres33_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1176 = {15'h0,io_in_bits_Pctrl_mulres33_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_172 = _T_1156 ? _T_1175 : _T_1176; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_226 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_172} : 34'h0; // @[PMDU.scala 1051:39 1081:30]
  wire [33:0] _GEN_247 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_226; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_260 = io_in_bits_Pctrl_isS1632 ? {{32'd0}, _T_1051} : _GEN_247; // @[PMDU.scala 1000:41 1023:30]
  wire [33:0] _GEN_278 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_260; // @[PMDU.scala 963:44]
  wire [33:0] adder34_3_1 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_278; // @[PMDU.scala 929:38]
  wire [14:0] _T_1135 = io_in_bits_Pctrl_mulres9_2[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1136 = {_T_1135,io_in_bits_Pctrl_mulres9_2[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1137 = {15'h0,io_in_bits_Pctrl_mulres9_2[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_168 = _T_1156 ? _T_1136 : _T_1137; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_221 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_168} : 34'h0; // @[PMDU.scala 1051:39 1081:30]
  wire [33:0] _GEN_242 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_221; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_255 = io_in_bits_Pctrl_isS1632 ? {{32'd0}, _T_1051} : _GEN_242; // @[PMDU.scala 1000:41 1023:30]
  wire [33:0] _GEN_277 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_255; // @[PMDU.scala 963:44]
  wire [33:0] adder34_3_0 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_277; // @[PMDU.scala 929:38]
  wire [70:0] _T_15 = {adder34_3_1,3'h0,adder34_3_0}; // @[Cat.scala 30:58]
  wire [1:0] _T_574 = _T_541 + _T_546; // @[PMDU.scala 911:46]
  wire [70:0] _GEN_69 = io_in_bits_Pctrl_isPMA_64ONLY ? {{69'd0}, _T_574} : _T_15; // @[PMDU.scala 731:15 902:50 911:27]
  wire [70:0] _GEN_77 = io_in_bits_Pctrl_isQ63_64ONLY ? _T_15 : _GEN_69; // @[PMDU.scala 731:15 886:50]
  wire [70:0] _GEN_83 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_15 : _GEN_77; // @[PMDU.scala 731:15 884:53]
  wire [70:0] _GEN_95 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_15 : _GEN_83; // @[PMDU.scala 731:15 836:50]
  wire [70:0] _GEN_107 = io_in_bits_Pctrl_isMul_8 ? _T_15 : _GEN_95; // @[PMDU.scala 731:15 779:45]
  wire [70:0] _GEN_119 = io_in_bits_Pctrl_isMul_16 ? _T_15 : _GEN_107; // @[PMDU.scala 731:15 735:40]
  wire [1:0] _T_1223 = {io_out_bits_DecodeOut_ctrl_fuOpType[0],1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1298 = _T_1266 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1272 = _T_467 ? io_in_bits_Pctrl_mulres65_0[31:0] : io_in_bits_Pctrl_mulres17_1[31:0]; // @[PMDU.scala 1133:23]
  wire [31:0] _T_1301 = _T_1272[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1302 = {_T_1301,_T_1272}; // @[Cat.scala 30:58]
  wire [63:0] _T_1303 = _T_1298 ^ _T_1302; // @[PMDU.scala 1139:50]
  wire [70:0] _GEN_207 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1303} : _GEN_119; // @[PMDU.scala 1126:40 1139:23]
  wire [70:0] _GEN_214 = io_in_bits_Pctrl_is3264 ? {{69'd0}, _T_1223} : _GEN_207; // @[PMDU.scala 1089:40 1101:23]
  wire [70:0] _GEN_232 = io_in_bits_Pctrl_is832 ? _GEN_119 : _GEN_214; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_249 = io_in_bits_Pctrl_isS1664 ? _GEN_119 : _GEN_232; // @[PMDU.scala 1046:41]
  wire [70:0] _GEN_267 = io_in_bits_Pctrl_isS1632 ? _GEN_119 : _GEN_249; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_284 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_119 : _GEN_267; // @[PMDU.scala 963:44]
  wire [70:0] adder68_3 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_119 : _GEN_284; // @[PMDU.scala 929:38]
  wire [70:0] _T_9 = _T_7 + adder68_3; // @[PMDU.scala 726:48]
  wire [14:0] _T_1181 = io_in_bits_Pctrl_mulres65_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1182 = {_T_1181,io_in_bits_Pctrl_mulres65_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1183 = {15'h0,io_in_bits_Pctrl_mulres65_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_173 = _T_1156 ? _T_1182 : _T_1183; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_227 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_173} : 34'h0; // @[PMDU.scala 1051:39 1082:30]
  wire [33:0] _GEN_248 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_227; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_266 = io_in_bits_Pctrl_isS1632 ? 34'h0 : _GEN_248; // @[PMDU.scala 1000:41]
  wire [33:0] _GEN_283 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_266; // @[PMDU.scala 963:44]
  wire [33:0] adder34_4_1 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_283; // @[PMDU.scala 929:38]
  wire [14:0] _T_1142 = io_in_bits_Pctrl_mulres9_3[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1143 = {_T_1142,io_in_bits_Pctrl_mulres9_3[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1144 = {15'h0,io_in_bits_Pctrl_mulres9_3[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_169 = _T_1156 ? _T_1143 : _T_1144; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_222 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_169} : 34'h0; // @[PMDU.scala 1051:39 1082:30]
  wire [33:0] _GEN_243 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_222; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_265 = io_in_bits_Pctrl_isS1632 ? 34'h0 : _GEN_243; // @[PMDU.scala 1000:41]
  wire [33:0] _GEN_282 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_265; // @[PMDU.scala 963:44]
  wire [33:0] adder34_4_0 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_282; // @[PMDU.scala 929:38]
  wire [70:0] _T_16 = {adder34_4_1,3'h0,adder34_4_0}; // @[Cat.scala 30:58]
  wire [31:0] _T_1276 = _T_467 ? 32'h0 : io_in_bits_Pctrl_mulres65_0[31:0]; // @[PMDU.scala 1135:23]
  wire [31:0] _T_1308 = _T_1276[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1309 = {_T_1308,_T_1276}; // @[Cat.scala 30:58]
  wire [63:0] _T_1310 = _T_1298 ^ _T_1309; // @[PMDU.scala 1140:50]
  wire [70:0] _GEN_208 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1310} : _T_16; // @[PMDU.scala 1126:40 1140:23 732:15]
  wire [70:0] _GEN_217 = io_in_bits_Pctrl_is3264 ? _T_16 : _GEN_208; // @[PMDU.scala 1089:40 732:15]
  wire [70:0] _GEN_234 = io_in_bits_Pctrl_is832 ? _T_16 : _GEN_217; // @[PMDU.scala 1051:39 732:15]
  wire [70:0] _GEN_251 = io_in_bits_Pctrl_isS1664 ? _T_16 : _GEN_234; // @[PMDU.scala 1046:41 732:15]
  wire [70:0] _GEN_268 = io_in_bits_Pctrl_isS1632 ? _T_16 : _GEN_251; // @[PMDU.scala 1000:41 732:15]
  wire [70:0] _GEN_285 = io_in_bits_Pctrl_isMSW_3216 ? _T_16 : _GEN_268; // @[PMDU.scala 732:15 963:44]
  wire [70:0] adder68_4 = io_in_bits_Pctrl_isMSW_3232 ? _T_16 : _GEN_285; // @[PMDU.scala 732:15 929:38]
  wire [70:0] tmp68 = _T_9 + adder68_4; // @[PMDU.scala 726:60]
  wire  _T_21 = io_out_bits_DecodeOut_ctrl_fuOpType[1:0] == 2'h1 | io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h9; // @[PMDU.scala 671:57]
  wire [15:0] _GEN_0 = _T_21 ? io_out_bits_DecodeOut_data_src2[31:16] : io_out_bits_DecodeOut_data_src2[15:0]; // @[PMDU.scala 687:23 689:29]
  wire [15:0] _GEN_1 = _T_21 ? io_out_bits_DecodeOut_data_src2[15:0] : io_out_bits_DecodeOut_data_src2[31:16]; // @[PMDU.scala 687:23 691:29]
  wire [15:0] _GEN_2 = _T_21 ? io_out_bits_DecodeOut_data_src2[63:48] : io_out_bits_DecodeOut_data_src2[47:32]; // @[PMDU.scala 687:23 689:29]
  wire [15:0] _GEN_3 = _T_21 ? io_out_bits_DecodeOut_data_src2[47:32] : io_out_bits_DecodeOut_data_src2[63:48]; // @[PMDU.scala 687:23 691:29]
  wire [63:0] _T_32 = {_GEN_3,_GEN_2,_GEN_1,_GEN_0}; // @[Cat.scala 30:58]
  wire  _T_34 = io_out_bits_DecodeOut_ctrl_fuOpType[1:0] == 2'h3; // @[PMDU.scala 672:44]
  wire [31:0] _T_48 = io_in_bits_Pctrl_mulres17_0[31:0]; // @[PMDU.scala 749:75]
  wire [16:0] _T_50 = _T_48[31:15]; // @[PMDU.scala 749:89]
  wire [31:0] _GEN_5 = _T_32[15:0] == 16'h8000 & io_out_bits_DecodeOut_data_src1[15:0] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_50}; // @[PMDU.scala 744:153 746:33 749:37]
  wire [31:0] _T_72 = io_in_bits_Pctrl_mulres17_1[31:0]; // @[PMDU.scala 751:75]
  wire [16:0] _T_74 = _T_72[31:15]; // @[PMDU.scala 751:89]
  wire [31:0] _GEN_7 = _T_32[31:16] == 16'h8000 & io_out_bits_DecodeOut_data_src1[31:16] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_74}; // @[PMDU.scala 744:153 746:33 751:37]
  wire [31:0] _T_96 = io_in_bits_Pctrl_mulres33_0[31:0]; // @[PMDU.scala 753:75]
  wire [16:0] _T_98 = _T_96[31:15]; // @[PMDU.scala 753:89]
  wire [31:0] _GEN_9 = _T_32[47:32] == 16'h8000 & io_out_bits_DecodeOut_data_src1[47:32] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_98}; // @[PMDU.scala 744:153 746:33 753:37]
  wire  _GEN_10 = _T_32[63:48] == 16'h8000 & io_out_bits_DecodeOut_data_src1[63:48] == 16'h8000 | (_T_32[47:32] == 16'h8000
     & io_out_bits_DecodeOut_data_src1[47:32] == 16'h8000 | (_T_32[31:16] == 16'h8000 & io_out_bits_DecodeOut_data_src1[
    31:16] == 16'h8000 | _T_32[15:0] == 16'h8000 & io_out_bits_DecodeOut_data_src1[15:0] == 16'h8000)); // @[PMDU.scala 744:153 745:59]
  wire [31:0] _GEN_11 = _T_32[63:48] == 16'h8000 & io_out_bits_DecodeOut_data_src1[63:48] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_1367}; // @[PMDU.scala 744:153 746:33 755:37]
  wire [63:0] _T_133 = {_GEN_11[15:0],_GEN_9[15:0],_GEN_7[15:0],_GEN_5[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_136 = {io_in_bits_Pctrl_mulres65_0[31:0],io_in_bits_Pctrl_mulres17_0[31:0]}; // @[Cat.scala 30:58]
  wire  _GEN_12 = _T_34 & _GEN_10; // @[PMDU.scala 705:35 738:39]
  wire [63:0] _GEN_13 = _T_34 ? _T_133 : _T_136; // @[PMDU.scala 738:39 739:36 764:36]
  wire [7:0] _GEN_14 = _T_21 ? io_out_bits_DecodeOut_data_src2[15:8] : io_out_bits_DecodeOut_data_src2[7:0]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_15 = _T_21 ? io_out_bits_DecodeOut_data_src2[7:0] : io_out_bits_DecodeOut_data_src2[15:8]; // @[PMDU.scala 687:23 691:29]
  wire [7:0] _GEN_16 = _T_21 ? io_out_bits_DecodeOut_data_src2[31:24] : io_out_bits_DecodeOut_data_src2[23:16]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_17 = _T_21 ? io_out_bits_DecodeOut_data_src2[23:16] : io_out_bits_DecodeOut_data_src2[31:24]; // @[PMDU.scala 687:23 691:29]
  wire [7:0] _GEN_18 = _T_21 ? io_out_bits_DecodeOut_data_src2[47:40] : io_out_bits_DecodeOut_data_src2[39:32]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_19 = _T_21 ? io_out_bits_DecodeOut_data_src2[39:32] : io_out_bits_DecodeOut_data_src2[47:40]; // @[PMDU.scala 687:23 691:29]
  wire [7:0] _GEN_20 = _T_21 ? io_out_bits_DecodeOut_data_src2[63:56] : io_out_bits_DecodeOut_data_src2[55:48]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_21 = _T_21 ? io_out_bits_DecodeOut_data_src2[55:48] : io_out_bits_DecodeOut_data_src2[63:56]; // @[PMDU.scala 687:23 691:29]
  wire [63:0] _T_164 = {_GEN_21,_GEN_20,_GEN_19,_GEN_18,_GEN_17,_GEN_16,_GEN_15,_GEN_14}; // @[Cat.scala 30:58]
  wire [15:0] _T_180 = io_in_bits_Pctrl_mulres9_0[15:0]; // @[PMDU.scala 793:74]
  wire [8:0] _T_182 = _T_180[15:7]; // @[PMDU.scala 793:87]
  wire [15:0] _GEN_23 = _T_164[7:0] == 8'h80 & io_out_bits_DecodeOut_data_src1[7:0] == 8'h80 ? 16'h7f : {{7'd0}, _T_182}
    ; // @[PMDU.scala 788:151 790:33 793:37]
  wire [15:0] _T_204 = io_in_bits_Pctrl_mulres9_1[15:0]; // @[PMDU.scala 795:74]
  wire [8:0] _T_206 = _T_204[15:7]; // @[PMDU.scala 795:87]
  wire [15:0] _GEN_25 = _T_164[15:8] == 8'h80 & io_out_bits_DecodeOut_data_src1[15:8] == 8'h80 ? 16'h7f : {{7'd0},
    _T_206}; // @[PMDU.scala 788:151 790:33 795:37]
  wire [15:0] _T_228 = io_in_bits_Pctrl_mulres9_2[15:0]; // @[PMDU.scala 797:74]
  wire [8:0] _T_230 = _T_228[15:7]; // @[PMDU.scala 797:87]
  wire [15:0] _GEN_27 = _T_164[23:16] == 8'h80 & io_out_bits_DecodeOut_data_src1[23:16] == 8'h80 ? 16'h7f : {{7'd0},
    _T_230}; // @[PMDU.scala 788:151 790:33 797:37]
  wire [15:0] _T_252 = io_in_bits_Pctrl_mulres9_3[15:0]; // @[PMDU.scala 799:74]
  wire [8:0] _T_254 = _T_252[15:7]; // @[PMDU.scala 799:87]
  wire [15:0] _GEN_29 = _T_164[31:24] == 8'h80 & io_out_bits_DecodeOut_data_src1[31:24] == 8'h80 ? 16'h7f : {{7'd0},
    _T_254}; // @[PMDU.scala 788:151 790:33 799:37]
  wire [15:0] _T_276 = io_in_bits_Pctrl_mulres17_0[15:0]; // @[PMDU.scala 801:75]
  wire [8:0] _T_278 = _T_276[15:7]; // @[PMDU.scala 801:88]
  wire [15:0] _GEN_31 = _T_164[39:32] == 8'h80 & io_out_bits_DecodeOut_data_src1[39:32] == 8'h80 ? 16'h7f : {{7'd0},
    _T_278}; // @[PMDU.scala 788:151 790:33 801:37]
  wire [15:0] _T_300 = io_in_bits_Pctrl_mulres17_1[15:0]; // @[PMDU.scala 803:75]
  wire [8:0] _T_302 = _T_300[15:7]; // @[PMDU.scala 803:88]
  wire [15:0] _GEN_33 = _T_164[47:40] == 8'h80 & io_out_bits_DecodeOut_data_src1[47:40] == 8'h80 ? 16'h7f : {{7'd0},
    _T_302}; // @[PMDU.scala 788:151 790:33 803:37]
  wire [15:0] _T_324 = io_in_bits_Pctrl_mulres33_0[15:0]; // @[PMDU.scala 805:75]
  wire [8:0] _T_326 = _T_324[15:7]; // @[PMDU.scala 805:88]
  wire  _GEN_34 = _T_164[55:48] == 8'h80 & io_out_bits_DecodeOut_data_src1[55:48] == 8'h80 | (_T_164[47:40] == 8'h80 &
    io_out_bits_DecodeOut_data_src1[47:40] == 8'h80 | (_T_164[39:32] == 8'h80 & io_out_bits_DecodeOut_data_src1[39:32]
     == 8'h80 | (_T_164[31:24] == 8'h80 & io_out_bits_DecodeOut_data_src1[31:24] == 8'h80 | (_T_164[23:16] == 8'h80 &
    io_out_bits_DecodeOut_data_src1[23:16] == 8'h80 | (_T_164[15:8] == 8'h80 & io_out_bits_DecodeOut_data_src1[15:8] == 8'h80
     | _T_164[7:0] == 8'h80 & io_out_bits_DecodeOut_data_src1[7:0] == 8'h80))))); // @[PMDU.scala 788:151 789:59]
  wire [15:0] _GEN_35 = _T_164[55:48] == 8'h80 & io_out_bits_DecodeOut_data_src1[55:48] == 8'h80 ? 16'h7f : {{7'd0},
    _T_326}; // @[PMDU.scala 788:151 790:33 805:37]
  wire [15:0] _T_348 = io_in_bits_Pctrl_mulres65_0[15:0]; // @[PMDU.scala 807:75]
  wire [8:0] _T_350 = _T_348[15:7]; // @[PMDU.scala 807:88]
  wire  _GEN_36 = _T_164[63:56] == 8'h80 & io_out_bits_DecodeOut_data_src1[63:56] == 8'h80 | _GEN_34; // @[PMDU.scala 788:151 789:59]
  wire [15:0] _GEN_37 = _T_164[63:56] == 8'h80 & io_out_bits_DecodeOut_data_src1[63:56] == 8'h80 ? 16'h7f : {{7'd0},
    _T_350}; // @[PMDU.scala 788:151 790:33 807:37]
  wire [63:0] _T_365 = {_GEN_37[7:0],_GEN_35[7:0],_GEN_33[7:0],_GEN_31[7:0],_GEN_29[7:0],_GEN_27[7:0],_GEN_25[7:0],
    _GEN_23[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_400 = {io_in_bits_Pctrl_mulres65_0[15:0],io_in_bits_Pctrl_mulres9_2[15:0],io_in_bits_Pctrl_mulres9_1[15
    :0],io_in_bits_Pctrl_mulres9_0[15:0]}; // @[Cat.scala 30:58]
  wire  _GEN_38 = _T_34 & _GEN_36; // @[PMDU.scala 705:35 782:39]
  wire [63:0] _GEN_39 = _T_34 ? _T_365 : _T_400; // @[PMDU.scala 782:39 783:36 816:36]
  wire [32:0] _T_445 = tmp68[32] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _GEN_304 = {{1'd0}, _T_445}; // @[PMDU.scala 870:63]
  wire [33:0] _T_447 = _GEN_304 ^ tmp68[33:0]; // @[PMDU.scala 870:63]
  wire  _T_449 = _T_447[32:31] != 2'h0; // @[PMDU.scala 870:92]
  wire [31:0] _GEN_44 = tmp68[32] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 872:65 873:36 875:37]
  wire  _GEN_45 = _T_447[32:31] != 2'h0 | _T_422; // @[PMDU.scala 870:100 871:59]
  wire [31:0] _GEN_46 = _T_447[32:31] != 2'h0 ? _GEN_44 : tmp68[31:0]; // @[PMDU.scala 870:100]
  wire  _GEN_47 = _T_467 ? _GEN_45 : _T_422; // @[PMDU.scala 869:53]
  wire [31:0] _GEN_48 = _T_467 ? _GEN_46 : tmp68[31:0]; // @[PMDU.scala 869:53]
  wire  _GEN_51 = _T_461 == 16'h8000 & _T_464 == 16'h8000 | _GEN_47; // @[PMDU.scala 851:77 852:55]
  wire [32:0] _T_497 = tmp68[69] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _GEN_305 = {{1'd0}, _T_497}; // @[PMDU.scala 870:63]
  wire [33:0] _T_499 = _GEN_305 ^ tmp68[70:37]; // @[PMDU.scala 870:63]
  wire  _T_501 = _T_499[32:31] != 2'h0; // @[PMDU.scala 870:92]
  wire [31:0] _GEN_53 = tmp68[69] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 872:65 873:36 875:37]
  wire  _GEN_54 = _T_499[32:31] != 2'h0 | _GEN_51; // @[PMDU.scala 870:100 871:59]
  wire [31:0] _GEN_55 = _T_499[32:31] != 2'h0 ? _GEN_53 : tmp68[68:37]; // @[PMDU.scala 870:100]
  wire  _GEN_56 = _T_467 ? _GEN_54 : _GEN_51; // @[PMDU.scala 869:53]
  wire [31:0] _GEN_57 = _T_467 ? _GEN_55 : tmp68[68:37]; // @[PMDU.scala 869:53]
  wire [63:0] _T_509 = {_GEN_57,_GEN_48}; // @[Cat.scala 30:58]
  wire [64:0] _T_519 = tmp68[64] ? 65'h1ffffffffffffffff : 65'h0; // @[Bitwise.scala 72:12]
  wire [70:0] _GEN_306 = {{6'd0}, _T_519}; // @[PMDU.scala 892:41]
  wire [70:0] _T_520 = _GEN_306 ^ tmp68; // @[PMDU.scala 892:41]
  wire  _T_522 = _T_520[64:63] != 2'h0; // @[PMDU.scala 892:56]
  wire [63:0] _GEN_58 = tmp68[64] ? 64'h8000000000000000 : 64'h7fffffffffffffff; // @[PMDU.scala 894:43 895:29 897:29]
  wire [63:0] _GEN_60 = _T_520[64:63] != 2'h0 ? _GEN_58 : tmp68[63:0]; // @[PMDU.scala 892:64]
  wire  _T_552 = ~(_T_924 & _T_467); // @[PMDU.scala 907:34]
  wire [65:0] _T_578 = tmp68[65] ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [70:0] _GEN_307 = {{5'd0}, _T_578}; // @[PMDU.scala 914:45]
  wire [70:0] _T_579 = _GEN_307 ^ tmp68; // @[PMDU.scala 914:45]
  wire  _T_581 = _T_579[65:63] != 3'h0; // @[PMDU.scala 914:59]
  wire [63:0] _GEN_61 = tmp68[65] ? 64'h8000000000000000 : 64'h7fffffffffffffff; // @[PMDU.scala 916:40 917:33 919:33]
  wire [63:0] _GEN_63 = _T_579[65:63] != 3'h0 ? _GEN_61 : tmp68[63:0]; // @[PMDU.scala 914:66]
  wire  _GEN_64 = _T_552 & _T_581; // @[PMDU.scala 913:33 705:35]
  wire [63:0] _GEN_65 = _T_552 ? _GEN_63 : tmp68[63:0]; // @[PMDU.scala 913:33]
  wire  _GEN_70 = io_in_bits_Pctrl_isPMA_64ONLY & _GEN_64; // @[PMDU.scala 705:35 902:50]
  wire [63:0] _GEN_71 = io_in_bits_Pctrl_isPMA_64ONLY ? _GEN_65 : 64'h0; // @[PMDU.scala 704:24 902:50 903:32]
  wire  _GEN_75 = io_in_bits_Pctrl_isQ63_64ONLY ? _T_522 : _GEN_70; // @[PMDU.scala 886:50]
  wire [63:0] _GEN_76 = io_in_bits_Pctrl_isQ63_64ONLY ? _GEN_60 : _GEN_71; // @[PMDU.scala 886:50 887:32]
  wire [63:0] _GEN_78 = io_in_bits_Pctrl_isMul_32_64ONLY ? io_in_bits_Pctrl_mulres65_0[63:0] : _GEN_76; // @[PMDU.scala 884:53 885:32]
  wire  _GEN_82 = io_in_bits_Pctrl_isMul_32_64ONLY ? 1'h0 : _GEN_75; // @[PMDU.scala 705:35 884:53]
  wire  _GEN_84 = io_in_bits_Pctrl_isQ15_64ONLY ? _GEN_56 : _GEN_82; // @[PMDU.scala 836:50]
  wire [63:0] _GEN_91 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_509 : _GEN_78; // @[PMDU.scala 836:50 837:32]
  wire  _GEN_96 = io_in_bits_Pctrl_isMul_8 ? _GEN_38 : _GEN_84; // @[PMDU.scala 779:45]
  wire [63:0] _GEN_97 = io_in_bits_Pctrl_isMul_8 ? _GEN_39 : _GEN_91; // @[PMDU.scala 779:45]
  wire  _GEN_108 = io_in_bits_Pctrl_isMul_16 ? _GEN_12 : _GEN_96; // @[PMDU.scala 735:40]
  wire [63:0] _GEN_109 = io_in_bits_Pctrl_isMul_16 ? _GEN_13 : _GEN_97; // @[PMDU.scala 735:40]
  wire  _T_612 = _T_694 & io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h0; // @[PMDU.scala 934:52]
  wire  _GEN_121 = _T_449 | _GEN_108; // @[PMDU.scala 945:96 946:55]
  wire  _GEN_123 = _T_803 & io_out_bits_DecodeOut_data_src2[31:0] == 32'h80000000 | _GEN_108; // @[PMDU.scala 954:147 955:55]
  wire [31:0] _GEN_124 = _T_803 & io_out_bits_DecodeOut_data_src2[31:0] == 32'h80000000 ? 32'h7fffffff : tmp68[31:0]; // @[PMDU.scala 954:147 956:29]
  wire  _GEN_125 = _T_697 ? _GEN_123 : _GEN_108; // @[PMDU.scala 953:32]
  wire [31:0] _GEN_126 = _T_697 ? _GEN_124 : tmp68[31:0]; // @[PMDU.scala 953:32]
  wire  _GEN_127 = _T_612 | _T_687 ? _GEN_121 : _GEN_125; // @[PMDU.scala 944:33]
  wire [31:0] _GEN_128 = _T_612 | _T_687 ? _GEN_46 : _GEN_126; // @[PMDU.scala 944:33]
  wire  _GEN_130 = _T_501 | _GEN_127; // @[PMDU.scala 945:96 946:55]
  wire  _GEN_132 = _T_880 & io_out_bits_DecodeOut_data_src2[63:32] == 32'h80000000 | _GEN_127; // @[PMDU.scala 954:147 955:55]
  wire [31:0] _GEN_133 = _T_880 & io_out_bits_DecodeOut_data_src2[63:32] == 32'h80000000 ? 32'h7fffffff : tmp68[68:37]; // @[PMDU.scala 954:147 956:29]
  wire  _GEN_134 = _T_697 ? _GEN_132 : _GEN_127; // @[PMDU.scala 953:32]
  wire [31:0] _GEN_135 = _T_697 ? _GEN_133 : tmp68[68:37]; // @[PMDU.scala 953:32]
  wire  _GEN_136 = _T_612 | _T_687 ? _GEN_130 : _GEN_134; // @[PMDU.scala 944:33]
  wire [31:0] _GEN_137 = _T_612 | _T_687 ? _GEN_55 : _GEN_135; // @[PMDU.scala 944:33]
  wire [63:0] _T_763 = {_GEN_137,_GEN_128}; // @[Cat.scala 30:58]
  wire  _T_768 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h3 | io_out_bits_DecodeOut_ctrl_fuOpType[6:5] == 2'h3; // @[PMDU.scala 967:54]
  wire  _GEN_138 = _T_847 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80000000 & _T_781 == 16'h8000 | _GEN_108; // @[PMDU.scala 975:127 976:51]
  wire  _GEN_141 = _T_449 | _GEN_138; // @[PMDU.scala 987:96 988:55]
  wire  _GEN_143 = _T_768 ? _GEN_141 : _GEN_138; // @[PMDU.scala 986:26]
  wire [31:0] _GEN_144 = _T_768 ? _GEN_46 : tmp68[31:0]; // @[PMDU.scala 986:26]
  wire  _GEN_145 = _T_847 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80000000 & _T_858 == 16'h8000 | _GEN_143; // @[PMDU.scala 975:127 976:51]
  wire  _GEN_148 = _T_501 | _GEN_145; // @[PMDU.scala 987:96 988:55]
  wire  _GEN_150 = _T_768 ? _GEN_148 : _GEN_145; // @[PMDU.scala 986:26]
  wire [31:0] _GEN_151 = _T_768 ? _GEN_55 : tmp68[68:37]; // @[PMDU.scala 986:26]
  wire [63:0] _T_918 = {_GEN_151,_GEN_144}; // @[Cat.scala 30:58]
  wire  _T_951 = io_out_bits_DecodeOut_ctrl_fuOpType[6:1] == 6'he; // @[PMDU.scala 1004:40]
  wire  _T_959 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h4 | _T_922 | _T_476; // @[PMDU.scala 1005:84]
  wire [31:0] _GEN_152 = _T_951 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80008000 &
    io_out_bits_DecodeOut_data_src2[31:0] == 32'h80008000 ? 32'h7fffffff : tmp68[31:0]; // @[PMDU.scala 1025:21 1026:211 1027:25]
  wire  _GEN_153 = _T_951 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80008000 & io_out_bits_DecodeOut_data_src2[31:0
    ] == 32'h80008000 | _GEN_108; // @[PMDU.scala 1026:211 1028:51]
  wire [33:0] _T_1008 = tmp68[33] ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1010 = _T_1008 ^ tmp68[33:0]; // @[PMDU.scala 1031:59]
  wire [31:0] _GEN_154 = tmp68[33] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 1033:61 1034:33 1036:33]
  wire  _GEN_155 = _T_1010[33:31] != 3'h0 | _GEN_153; // @[PMDU.scala 1031:96 1032:55]
  wire [31:0] _GEN_156 = _T_1010[33:31] != 3'h0 ? _GEN_154 : _GEN_152; // @[PMDU.scala 1031:96]
  wire  _GEN_157 = _T_959 ? _GEN_155 : _GEN_153; // @[PMDU.scala 1030:33]
  wire [31:0] _GEN_158 = _T_959 ? _GEN_156 : _GEN_152; // @[PMDU.scala 1030:33]
  wire [31:0] _GEN_159 = _T_951 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80008000 &
    io_out_bits_DecodeOut_data_src2[63:32] == 32'h80008000 ? 32'h7fffffff : tmp68[68:37]; // @[PMDU.scala 1025:21 1026:211 1027:25]
  wire  _GEN_160 = _T_951 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80008000 & io_out_bits_DecodeOut_data_src2[63:
    32] == 32'h80008000 | _GEN_157; // @[PMDU.scala 1026:211 1028:51]
  wire [33:0] _T_1075 = tmp68[70] ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1077 = _T_1075 ^ tmp68[70:37]; // @[PMDU.scala 1031:59]
  wire [31:0] _GEN_161 = tmp68[70] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 1033:61 1034:33 1036:33]
  wire  _GEN_162 = _T_1077[33:31] != 3'h0 | _GEN_160; // @[PMDU.scala 1031:96 1032:55]
  wire [31:0] _GEN_163 = _T_1077[33:31] != 3'h0 ? _GEN_161 : _GEN_159; // @[PMDU.scala 1031:96]
  wire  _GEN_164 = _T_959 ? _GEN_162 : _GEN_160; // @[PMDU.scala 1030:33]
  wire [31:0] _GEN_165 = _T_959 ? _GEN_163 : _GEN_159; // @[PMDU.scala 1030:33]
  wire [63:0] _T_1096 = {_GEN_165,_GEN_158}; // @[Cat.scala 30:58]
  wire [63:0] _T_1195 = {tmp68[68:37],tmp68[31:0]}; // @[Cat.scala 30:58]
  wire  _GEN_178 = _T_581 | _GEN_108; // @[PMDU.scala 1105:68 1106:55]
  wire  _GEN_180 = ~io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65:64] != 2'h0 | _GEN_108; // @[PMDU.scala 1117:61 1118:55]
  wire [63:0] _GEN_181 = ~io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65:64] != 2'h0 ? 64'hffffffffffffffff : tmp68[
    63:0]; // @[PMDU.scala 1117:61 1119:29]
  wire  _GEN_182 = io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65] | _GEN_180; // @[PMDU.scala 1114:52 1115:55]
  wire [63:0] _GEN_183 = io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65] ? 64'h0 : _GEN_181; // @[PMDU.scala 1114:52 1116:29]
  wire  _GEN_184 = _T_1198 ? _GEN_178 : _GEN_182; // @[PMDU.scala 1104:31]
  wire [63:0] _GEN_185 = _T_1198 ? _GEN_63 : _GEN_183; // @[PMDU.scala 1104:31]
  wire  _GEN_186 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _GEN_184 : _GEN_108; // @[PMDU.scala 1103:29]
  wire [63:0] _GEN_187 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _GEN_185 : tmp68[63:0]; // @[PMDU.scala 1103:29]
  wire  _GEN_188 = _T_1354 == 16'h8000 & _T_1357 == 16'h8000 | _GEN_108; // @[PMDU.scala 1161:70 1162:47]
  wire [31:0] _T_1387 = tmp68[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1388 = {_T_1387,tmp68[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1391 = tmp68[32] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [70:0] _GEN_313 = {{38'd0}, _T_1391}; // @[PMDU.scala 1172:41]
  wire [70:0] _T_1392 = _GEN_313 ^ tmp68; // @[PMDU.scala 1172:41]
  wire [63:0] _GEN_190 = tmp68[32] ? 64'hffffffff80000000 : 64'h7fffffff; // @[PMDU.scala 1174:43 1175:29 1177:29]
  wire  _GEN_191 = _T_1392[32:31] != 2'h0 | _GEN_188; // @[PMDU.scala 1172:64 1173:51]
  wire [63:0] _GEN_192 = _T_1392[32:31] != 2'h0 ? _GEN_190 : _T_1388; // @[PMDU.scala 1171:21 1172:64]
  wire [63:0] _GEN_193 = _T_686 ? _GEN_192 : _GEN_189; // @[PMDU.scala 1170:30]
  wire  _GEN_194 = _T_686 ? _GEN_191 : _GEN_188; // @[PMDU.scala 1170:30]
  wire [63:0] _T_1431 = io_out_bits_DecodeOut_ctrl_fuOpType[4] ? tmp68[63:0] : _T_1388; // @[PMDU.scala 1189:16]
  wire [63:0] _GEN_198 = io_in_bits_Pctrl_isC31 ? _T_1431 : _GEN_109; // @[PMDU.scala 1183:39 1184:28]
  wire  _GEN_199 = io_in_bits_Pctrl_isQ15orQ31 ? _GEN_194 : _GEN_108; // @[PMDU.scala 1149:44]
  wire [63:0] _GEN_202 = io_in_bits_Pctrl_isQ15orQ31 ? _GEN_193 : _GEN_198; // @[PMDU.scala 1149:44 1150:28]
  wire [63:0] _GEN_209 = io_in_bits_Pctrl_is1664 ? tmp68[63:0] : _GEN_202; // @[PMDU.scala 1126:40 1130:28]
  wire  _GEN_210 = io_in_bits_Pctrl_is1664 ? _GEN_108 : _GEN_199; // @[PMDU.scala 1126:40]
  wire  _GEN_215 = io_in_bits_Pctrl_is3264 ? _GEN_186 : _GEN_210; // @[PMDU.scala 1089:40]
  wire [63:0] _GEN_216 = io_in_bits_Pctrl_is3264 ? _GEN_187 : _GEN_209; // @[PMDU.scala 1089:40 1093:28]
  wire [63:0] _GEN_228 = io_in_bits_Pctrl_is832 ? _T_1195 : _GEN_216; // @[PMDU.scala 1051:39 1053:28]
  wire  _GEN_233 = io_in_bits_Pctrl_is832 ? _GEN_108 : _GEN_215; // @[PMDU.scala 1051:39]
  wire [63:0] _GEN_238 = io_in_bits_Pctrl_isS1664 ? tmp68[63:0] : _GEN_228; // @[PMDU.scala 1046:41 1050:28]
  wire  _GEN_250 = io_in_bits_Pctrl_isS1664 ? _GEN_108 : _GEN_233; // @[PMDU.scala 1046:41]
  wire  _GEN_256 = io_in_bits_Pctrl_isS1632 ? _GEN_164 : _GEN_250; // @[PMDU.scala 1000:41]
  wire [63:0] _GEN_261 = io_in_bits_Pctrl_isS1632 ? _T_1096 : _GEN_238; // @[PMDU.scala 1000:41 1006:28]
  wire  _GEN_269 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_150 : _GEN_256; // @[PMDU.scala 963:44]
  wire [63:0] _GEN_276 = io_in_bits_Pctrl_isMSW_3216 ? _T_918 : _GEN_261; // @[PMDU.scala 963:44 964:28]
  assign io_in_ready = _T | ~io_in_valid; // @[PMDU.scala 701:35]
  assign io_out_valid = io_in_valid; // @[PMDU.scala 700:18]
  assign io_out_bits_result = io_in_bits_Pctrl_isMSW_3232 ? _T_763 : _GEN_276; // @[PMDU.scala 929:38 930:28]
  assign io_out_bits_DecodeOut_cf_pc = io_in_bits_DecodeIn_cf_pc; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_cf_runahead_checkpoint_id = io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_ctrl_fuOpType = io_in_bits_DecodeIn_ctrl_fuOpType; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_ctrl_rfWen = io_in_bits_DecodeIn_ctrl_rfWen; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_ctrl_rfDest = io_in_bits_DecodeIn_ctrl_rfDest; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_data_src1 = io_in_bits_DecodeIn_data_src1; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_data_src2 = io_in_bits_DecodeIn_data_src2; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_data_src3 = io_in_bits_DecodeIn_data_src3; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_pext_OV = io_in_bits_Pctrl_isMSW_3232 ? _GEN_136 : _GEN_269; // @[PMDU.scala 929:38]
  assign io_out_bits_DecodeOut_InstNo = io_in_bits_DecodeIn_InstNo; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_InstFlag = io_in_bits_DecodeIn_InstFlag; // @[PMDU.scala 703:27]
  assign io_FirstStageFire = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
endmodule
module PALU_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [38:0] io_in_bits_DecodeIn_cf_pc,
  input  [63:0] io_in_bits_DecodeIn_cf_runahead_checkpoint_id,
  input  [6:0]  io_in_bits_DecodeIn_ctrl_fuOpType,
  input  [2:0]  io_in_bits_DecodeIn_ctrl_funct3,
  input         io_in_bits_DecodeIn_ctrl_func24,
  input         io_in_bits_DecodeIn_ctrl_rfWen,
  input  [4:0]  io_in_bits_DecodeIn_ctrl_rfDest,
  input  [63:0] io_in_bits_DecodeIn_data_src1,
  input  [63:0] io_in_bits_DecodeIn_data_src2,
  input  [63:0] io_in_bits_DecodeIn_data_src3,
  input  [4:0]  io_in_bits_DecodeIn_InstNo,
  input         io_in_bits_DecodeIn_InstFlag,
  input         io_in_bits_Pctrl_isAdd_64,
  input         io_in_bits_Pctrl_isAdd_32,
  input         io_in_bits_Pctrl_isAdd_16,
  input         io_in_bits_Pctrl_isAdd_8,
  input         io_in_bits_Pctrl_isAdd_Q15,
  input         io_in_bits_Pctrl_isAdd_Q31,
  input         io_in_bits_Pctrl_isAdd_C31,
  input         io_in_bits_Pctrl_isAve,
  input         io_in_bits_Pctrl_isSub_64,
  input         io_in_bits_Pctrl_isSub_32,
  input         io_in_bits_Pctrl_isSub_16,
  input         io_in_bits_Pctrl_isSub_8,
  input         io_in_bits_Pctrl_isSub_Q15,
  input         io_in_bits_Pctrl_isSub_Q31,
  input         io_in_bits_Pctrl_isSub_C31,
  input         io_in_bits_Pctrl_isCras_16,
  input         io_in_bits_Pctrl_isCrsa_16,
  input         io_in_bits_Pctrl_isCras_32,
  input         io_in_bits_Pctrl_isCrsa_32,
  input         io_in_bits_Pctrl_isStas_16,
  input         io_in_bits_Pctrl_isStsa_16,
  input         io_in_bits_Pctrl_isStas_32,
  input         io_in_bits_Pctrl_isStsa_32,
  input         io_in_bits_Pctrl_isComp_16,
  input         io_in_bits_Pctrl_isComp_8,
  input         io_in_bits_Pctrl_isCompare,
  input         io_in_bits_Pctrl_isMaxMin_16,
  input         io_in_bits_Pctrl_isMaxMin_8,
  input         io_in_bits_Pctrl_isMaxMin_XLEN,
  input         io_in_bits_Pctrl_isMaxMin_32,
  input         io_in_bits_Pctrl_isMaxMin,
  input         io_in_bits_Pctrl_isPbs,
  input         io_in_bits_Pctrl_isRs_16,
  input         io_in_bits_Pctrl_isLs_16,
  input         io_in_bits_Pctrl_isLR_16,
  input         io_in_bits_Pctrl_isRs_8,
  input         io_in_bits_Pctrl_isLs_8,
  input         io_in_bits_Pctrl_isLR_8,
  input         io_in_bits_Pctrl_isRs_32,
  input         io_in_bits_Pctrl_isLs_32,
  input         io_in_bits_Pctrl_isLR_32,
  input         io_in_bits_Pctrl_isLR_Q31,
  input         io_in_bits_Pctrl_isLs_Q31,
  input         io_in_bits_Pctrl_isRs_XLEN,
  input         io_in_bits_Pctrl_isSRAIWU,
  input         io_in_bits_Pctrl_isFSRW,
  input         io_in_bits_Pctrl_isWext,
  input         io_in_bits_Pctrl_isShifter,
  input         io_in_bits_Pctrl_isClip_16,
  input         io_in_bits_Pctrl_isClip_8,
  input         io_in_bits_Pctrl_isclip_32,
  input         io_in_bits_Pctrl_isClip,
  input         io_in_bits_Pctrl_isSat_16,
  input         io_in_bits_Pctrl_isSat_8,
  input         io_in_bits_Pctrl_isSat_32,
  input         io_in_bits_Pctrl_isSat_W,
  input         io_in_bits_Pctrl_isSat,
  input         io_in_bits_Pctrl_isCnt_16,
  input         io_in_bits_Pctrl_isCnt_8,
  input         io_in_bits_Pctrl_isCnt_32,
  input         io_in_bits_Pctrl_isCnt,
  input         io_in_bits_Pctrl_isSwap_16,
  input         io_in_bits_Pctrl_isSwap_8,
  input         io_in_bits_Pctrl_isSwap,
  input         io_in_bits_Pctrl_isUnpack,
  input         io_in_bits_Pctrl_isBitrev,
  input         io_in_bits_Pctrl_isCmix,
  input         io_in_bits_Pctrl_isInsertb,
  input         io_in_bits_Pctrl_isPackbb,
  input         io_in_bits_Pctrl_isPackbt,
  input         io_in_bits_Pctrl_isPacktb,
  input         io_in_bits_Pctrl_isPacktt,
  input         io_in_bits_Pctrl_isPack,
  input  [7:0]  io_in_bits_Pctrl_isSub,
  input         io_in_bits_Pctrl_isAdder,
  input         io_in_bits_Pctrl_SrcSigned,
  input         io_in_bits_Pctrl_Saturating,
  input         io_in_bits_Pctrl_Translation,
  input         io_in_bits_Pctrl_LessEqual,
  input         io_in_bits_Pctrl_LessThan,
  input  [79:0] io_in_bits_Pctrl_adderRes_ori,
  input  [63:0] io_in_bits_Pctrl_adderRes,
  input  [79:0] io_in_bits_Pctrl_adderRes_ori_drophighestbit,
  input         io_in_bits_Pctrl_Round,
  input         io_in_bits_Pctrl_ShiftSigned,
  input         io_in_bits_Pctrl_Arithmetic,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_result,
  output [38:0] io_out_bits_DecodeOut_cf_pc,
  output [63:0] io_out_bits_DecodeOut_cf_runahead_checkpoint_id,
  output        io_out_bits_DecodeOut_ctrl_rfWen,
  output [4:0]  io_out_bits_DecodeOut_ctrl_rfDest,
  output        io_out_bits_DecodeOut_pext_OV,
  output [4:0]  io_out_bits_DecodeOut_InstNo,
  output        io_out_bits_DecodeOut_InstFlag
);
  wire  _T_1 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15; // @[PALU.scala 186:43]
  wire  _T_15 = ~io_in_bits_DecodeIn_ctrl_fuOpType[3]; // @[PALU.scala 186:55]
  wire  _T_16 = io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15 ? ~io_in_bits_DecodeIn_ctrl_fuOpType[3] :
    io_in_bits_Pctrl_SrcSigned; // @[PALU.scala 186:33]
  wire  _GEN_7 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[17] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[15] :
    io_in_bits_Pctrl_adderRes_ori[16]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_0 = io_in_bits_Pctrl_adderRes_ori[17] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_1 = _GEN_7 ? _GEN_0 : io_in_bits_Pctrl_adderRes_ori[15:0]; // @[PALU.scala 123:21 126:33]
  wire [15:0] _GEN_3 = io_in_bits_Pctrl_isSub[0] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_5 = _GEN_7 ? _GEN_3 : io_in_bits_Pctrl_adderRes_ori[15:0]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_8 = _T_16 ? _GEN_1 : _GEN_5; // @[PALU.scala 124:28]
  wire  _GEN_17 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[35] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[33] :
    io_in_bits_Pctrl_adderRes_ori[34]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_10 = io_in_bits_Pctrl_adderRes_ori[35] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_11 = _GEN_17 ? _GEN_10 : io_in_bits_Pctrl_adderRes_ori[33:18]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_12 = _GEN_17 | _GEN_7; // @[PALU.scala 126:33 132:24]
  wire [15:0] _GEN_13 = io_in_bits_Pctrl_isSub[1] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_15 = _GEN_17 ? _GEN_13 : io_in_bits_Pctrl_adderRes_ori[33:18]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_18 = _T_16 ? _GEN_11 : _GEN_15; // @[PALU.scala 124:28]
  wire  _GEN_19 = _T_16 ? _GEN_12 : _GEN_12; // @[PALU.scala 124:28]
  wire  _GEN_27 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[53] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[51] :
    io_in_bits_Pctrl_adderRes_ori[52]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_20 = io_in_bits_Pctrl_adderRes_ori[53] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_21 = _GEN_27 ? _GEN_20 : io_in_bits_Pctrl_adderRes_ori[51:36]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_22 = _GEN_27 | _GEN_19; // @[PALU.scala 126:33 132:24]
  wire [15:0] _GEN_23 = io_in_bits_Pctrl_isSub[2] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_25 = _GEN_27 ? _GEN_23 : io_in_bits_Pctrl_adderRes_ori[51:36]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_28 = _T_16 ? _GEN_21 : _GEN_25; // @[PALU.scala 124:28]
  wire  _GEN_29 = _T_16 ? _GEN_22 : _GEN_22; // @[PALU.scala 124:28]
  wire  _GEN_37 = _T_16 ? io_in_bits_Pctrl_adderRes_ori[71] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[69] :
    io_in_bits_Pctrl_adderRes_ori[70]; // @[PALU.scala 124:28 125:21 135:21]
  wire [15:0] _GEN_30 = io_in_bits_Pctrl_adderRes_ori[71] ? 16'h8000 : 16'h7fff; // @[PALU.scala 127:66 128:33 130:33]
  wire [15:0] _GEN_31 = _GEN_37 ? _GEN_30 : io_in_bits_Pctrl_adderRes_ori[69:54]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_32 = _GEN_37 | _GEN_29; // @[PALU.scala 126:33 132:24]
  wire [15:0] _GEN_33 = io_in_bits_Pctrl_isSub[3] ? 16'h0 : 16'hffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [15:0] _GEN_35 = _GEN_37 ? _GEN_33 : io_in_bits_Pctrl_adderRes_ori[69:54]; // @[PALU.scala 123:21 136:33]
  wire [15:0] _GEN_38 = _T_16 ? _GEN_31 : _GEN_35; // @[PALU.scala 124:28]
  wire  _GEN_39 = _T_16 ? _GEN_32 : _GEN_32; // @[PALU.scala 124:28]
  wire [64:0] _T_80 = {_GEN_39,_GEN_38,_GEN_28,_GEN_18,_GEN_8}; // @[Cat.scala 30:58]
  wire [47:0] _T_85 = _T_80[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_86 = {_T_85,_T_80[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_88 = _T_12 ? _T_86 : _T_80[63:0]; // @[PALU.scala 188:34]
  wire [63:0] _T_101 = {io_in_bits_Pctrl_adderRes_ori[70:55],io_in_bits_Pctrl_adderRes_ori[52:37],
    io_in_bits_Pctrl_adderRes_ori[34:19],io_in_bits_Pctrl_adderRes_ori[16:1]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_40 = io_in_bits_Pctrl_Translation ? _T_101 : io_in_bits_Pctrl_adderRes; // @[PALU.scala 190:32 191:28]
  wire [63:0] _GEN_41 = io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15 ? _T_88 :
    _GEN_40; // @[PALU.scala 185:49 188:28]
  wire  _GEN_42 = (io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q15 | io_in_bits_Pctrl_isSub_Q15) & _T_80[64]; // @[PALU.scala 185:49 189:21]
  wire  _GEN_50 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[9] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[7] : io_in_bits_Pctrl_adderRes_ori[8]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_43 = io_in_bits_Pctrl_adderRes_ori[9] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_44 = _GEN_50 ? _GEN_43 : io_in_bits_Pctrl_adderRes_ori[7:0]; // @[PALU.scala 123:21 126:33]
  wire [7:0] _GEN_46 = io_in_bits_Pctrl_isSub[0] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_48 = _GEN_50 ? _GEN_46 : io_in_bits_Pctrl_adderRes_ori[7:0]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_51 = io_in_bits_Pctrl_SrcSigned ? _GEN_44 : _GEN_48; // @[PALU.scala 124:28]
  wire  _GEN_60 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[19] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[17] : io_in_bits_Pctrl_adderRes_ori[18]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_53 = io_in_bits_Pctrl_adderRes_ori[19] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_54 = _GEN_60 ? _GEN_53 : io_in_bits_Pctrl_adderRes_ori[17:10]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_55 = _GEN_60 | _GEN_50; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_56 = io_in_bits_Pctrl_isSub[1] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_58 = _GEN_60 ? _GEN_56 : io_in_bits_Pctrl_adderRes_ori[17:10]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_61 = io_in_bits_Pctrl_SrcSigned ? _GEN_54 : _GEN_58; // @[PALU.scala 124:28]
  wire  _GEN_62 = io_in_bits_Pctrl_SrcSigned ? _GEN_55 : _GEN_55; // @[PALU.scala 124:28]
  wire  _GEN_70 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[29] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[27] : io_in_bits_Pctrl_adderRes_ori[28]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_63 = io_in_bits_Pctrl_adderRes_ori[29] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_64 = _GEN_70 ? _GEN_63 : io_in_bits_Pctrl_adderRes_ori[27:20]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_65 = _GEN_70 | _GEN_62; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_66 = io_in_bits_Pctrl_isSub[2] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_68 = _GEN_70 ? _GEN_66 : io_in_bits_Pctrl_adderRes_ori[27:20]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_71 = io_in_bits_Pctrl_SrcSigned ? _GEN_64 : _GEN_68; // @[PALU.scala 124:28]
  wire  _GEN_72 = io_in_bits_Pctrl_SrcSigned ? _GEN_65 : _GEN_65; // @[PALU.scala 124:28]
  wire  _GEN_80 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[39] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[37] : io_in_bits_Pctrl_adderRes_ori[38]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_73 = io_in_bits_Pctrl_adderRes_ori[39] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_74 = _GEN_80 ? _GEN_73 : io_in_bits_Pctrl_adderRes_ori[37:30]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_75 = _GEN_80 | _GEN_72; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_76 = io_in_bits_Pctrl_isSub[3] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_78 = _GEN_80 ? _GEN_76 : io_in_bits_Pctrl_adderRes_ori[37:30]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_81 = io_in_bits_Pctrl_SrcSigned ? _GEN_74 : _GEN_78; // @[PALU.scala 124:28]
  wire  _GEN_82 = io_in_bits_Pctrl_SrcSigned ? _GEN_75 : _GEN_75; // @[PALU.scala 124:28]
  wire  _GEN_90 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[49] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[47] : io_in_bits_Pctrl_adderRes_ori[48]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_83 = io_in_bits_Pctrl_adderRes_ori[49] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_84 = _GEN_90 ? _GEN_83 : io_in_bits_Pctrl_adderRes_ori[47:40]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_85 = _GEN_90 | _GEN_82; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_86 = io_in_bits_Pctrl_isSub[4] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_88 = _GEN_90 ? _GEN_86 : io_in_bits_Pctrl_adderRes_ori[47:40]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_91 = io_in_bits_Pctrl_SrcSigned ? _GEN_84 : _GEN_88; // @[PALU.scala 124:28]
  wire  _GEN_92 = io_in_bits_Pctrl_SrcSigned ? _GEN_85 : _GEN_85; // @[PALU.scala 124:28]
  wire  _GEN_100 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[59] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[57] : io_in_bits_Pctrl_adderRes_ori[58]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_93 = io_in_bits_Pctrl_adderRes_ori[59] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_94 = _GEN_100 ? _GEN_93 : io_in_bits_Pctrl_adderRes_ori[57:50]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_95 = _GEN_100 | _GEN_92; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_96 = io_in_bits_Pctrl_isSub[5] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_98 = _GEN_100 ? _GEN_96 : io_in_bits_Pctrl_adderRes_ori[57:50]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_101 = io_in_bits_Pctrl_SrcSigned ? _GEN_94 : _GEN_98; // @[PALU.scala 124:28]
  wire  _GEN_102 = io_in_bits_Pctrl_SrcSigned ? _GEN_95 : _GEN_95; // @[PALU.scala 124:28]
  wire  _GEN_110 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[69] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[67] : io_in_bits_Pctrl_adderRes_ori[68]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_103 = io_in_bits_Pctrl_adderRes_ori[69] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_104 = _GEN_110 ? _GEN_103 : io_in_bits_Pctrl_adderRes_ori[67:60]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_105 = _GEN_110 | _GEN_102; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_106 = io_in_bits_Pctrl_isSub[6] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_108 = _GEN_110 ? _GEN_106 : io_in_bits_Pctrl_adderRes_ori[67:60]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_111 = io_in_bits_Pctrl_SrcSigned ? _GEN_104 : _GEN_108; // @[PALU.scala 124:28]
  wire  _GEN_112 = io_in_bits_Pctrl_SrcSigned ? _GEN_105 : _GEN_105; // @[PALU.scala 124:28]
  wire  _GEN_120 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[79] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[77] : io_in_bits_Pctrl_adderRes_ori[78]; // @[PALU.scala 124:28 125:21 135:21]
  wire [7:0] _GEN_113 = io_in_bits_Pctrl_adderRes_ori[79] ? 8'h80 : 8'h7f; // @[PALU.scala 127:66 128:33 130:33]
  wire [7:0] _GEN_114 = _GEN_120 ? _GEN_113 : io_in_bits_Pctrl_adderRes_ori[77:70]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_115 = _GEN_120 | _GEN_112; // @[PALU.scala 126:33 132:24]
  wire [7:0] _GEN_116 = io_in_bits_Pctrl_isSub[7] ? 8'h0 : 8'hff; // @[PALU.scala 137:35 138:33 141:33]
  wire [7:0] _GEN_118 = _GEN_120 ? _GEN_116 : io_in_bits_Pctrl_adderRes_ori[77:70]; // @[PALU.scala 123:21 136:33]
  wire [7:0] _GEN_121 = io_in_bits_Pctrl_SrcSigned ? _GEN_114 : _GEN_118; // @[PALU.scala 124:28]
  wire  _GEN_122 = io_in_bits_Pctrl_SrcSigned ? _GEN_115 : _GEN_115; // @[PALU.scala 124:28]
  wire [64:0] _T_230 = {_GEN_122,_GEN_121,_GEN_111,_GEN_101,_GEN_91,_GEN_81,_GEN_71,_GEN_61,_GEN_51}; // @[Cat.scala 30:58]
  wire [63:0] _T_256 = {io_in_bits_Pctrl_adderRes_ori[78:71],io_in_bits_Pctrl_adderRes_ori[68:61],
    io_in_bits_Pctrl_adderRes_ori[58:51],io_in_bits_Pctrl_adderRes_ori[48:41],io_in_bits_Pctrl_adderRes_ori[38:31],
    io_in_bits_Pctrl_adderRes_ori[28:21],io_in_bits_Pctrl_adderRes_ori[18:11],io_in_bits_Pctrl_adderRes_ori[8:1]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_123 = io_in_bits_Pctrl_Translation ? _T_256 : io_in_bits_Pctrl_adderRes; // @[PALU.scala 198:32 199:28]
  wire [63:0] _GEN_124 = io_in_bits_Pctrl_Saturating ? _T_230[63:0] : _GEN_123; // @[PALU.scala 194:25 196:28]
  wire  _GEN_125 = io_in_bits_Pctrl_Saturating & _T_230[64]; // @[PALU.scala 194:25 197:21]
  wire  _T_266 = io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31; // @[PALU.scala 203:44]
  wire  _T_270 = io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31 ? _T_15 : io_in_bits_Pctrl_SrcSigned; // @[PALU.scala 203:33]
  wire  _GEN_133 = _T_270 ? io_in_bits_Pctrl_adderRes_ori[33] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[31] :
    io_in_bits_Pctrl_adderRes_ori[32]; // @[PALU.scala 124:28 125:21 135:21]
  wire [31:0] _GEN_126 = io_in_bits_Pctrl_adderRes_ori[33] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 127:66 128:33 130:33]
  wire [31:0] _GEN_127 = _GEN_133 ? _GEN_126 : io_in_bits_Pctrl_adderRes_ori[31:0]; // @[PALU.scala 123:21 126:33]
  wire [31:0] _GEN_129 = io_in_bits_Pctrl_isSub[0] ? 32'h0 : 32'hffffffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [31:0] _GEN_131 = _GEN_133 ? _GEN_129 : io_in_bits_Pctrl_adderRes_ori[31:0]; // @[PALU.scala 123:21 136:33]
  wire [31:0] _GEN_134 = _T_270 ? _GEN_127 : _GEN_131; // @[PALU.scala 124:28]
  wire  _GEN_143 = _T_270 ? io_in_bits_Pctrl_adderRes_ori[67] ^ io_in_bits_Pctrl_adderRes_ori_drophighestbit[65] :
    io_in_bits_Pctrl_adderRes_ori[66]; // @[PALU.scala 124:28 125:21 135:21]
  wire [31:0] _GEN_136 = io_in_bits_Pctrl_adderRes_ori[67] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 127:66 128:33 130:33]
  wire [31:0] _GEN_137 = _GEN_143 ? _GEN_136 : io_in_bits_Pctrl_adderRes_ori[65:34]; // @[PALU.scala 123:21 126:33]
  wire  _GEN_138 = _GEN_143 | _GEN_133; // @[PALU.scala 126:33 132:24]
  wire [31:0] _GEN_139 = io_in_bits_Pctrl_isSub[1] ? 32'h0 : 32'hffffffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [31:0] _GEN_141 = _GEN_143 ? _GEN_139 : io_in_bits_Pctrl_adderRes_ori[65:34]; // @[PALU.scala 123:21 136:33]
  wire [31:0] _GEN_144 = _T_270 ? _GEN_137 : _GEN_141; // @[PALU.scala 124:28]
  wire  _GEN_145 = _T_270 ? _GEN_138 : _GEN_138; // @[PALU.scala 124:28]
  wire [64:0] _T_302 = {_GEN_145,_GEN_144,_GEN_134}; // @[Cat.scala 30:58]
  wire [31:0] _T_307 = _T_302[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_308 = {_T_307,_T_302[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_310 = _T_266 ? _T_308 : _T_302[63:0]; // @[PALU.scala 205:34]
  wire [63:0] _T_317 = {io_in_bits_Pctrl_adderRes_ori[66:35],io_in_bits_Pctrl_adderRes_ori[32:1]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_146 = io_in_bits_Pctrl_Translation ? _T_317 : io_in_bits_Pctrl_adderRes; // @[PALU.scala 207:32 208:28]
  wire [63:0] _GEN_147 = io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31 ? _T_310
     : _GEN_146; // @[PALU.scala 202:49 205:28]
  wire  _GEN_148 = (io_in_bits_Pctrl_Saturating | io_in_bits_Pctrl_isAdd_Q31 | io_in_bits_Pctrl_isSub_Q31) & _T_302[64]; // @[PALU.scala 202:49 206:21]
  wire  _GEN_156 = io_in_bits_Pctrl_SrcSigned ? io_in_bits_Pctrl_adderRes_ori[65] ^
    io_in_bits_Pctrl_adderRes_ori_drophighestbit[63] : io_in_bits_Pctrl_adderRes_ori[64]; // @[PALU.scala 124:28 125:21 135:21]
  wire [63:0] _GEN_149 = io_in_bits_Pctrl_adderRes_ori[65] ? 64'h8000000000000000 : 64'h7fffffffffffffff; // @[PALU.scala 127:66 128:33 130:33]
  wire [63:0] _GEN_150 = _GEN_156 ? _GEN_149 : io_in_bits_Pctrl_adderRes_ori[63:0]; // @[PALU.scala 123:21 126:33]
  wire [63:0] _GEN_152 = io_in_bits_Pctrl_isSub[0] ? 64'h0 : 64'hffffffffffffffff; // @[PALU.scala 137:35 138:33 141:33]
  wire [63:0] _GEN_154 = _GEN_156 ? _GEN_152 : io_in_bits_Pctrl_adderRes_ori[63:0]; // @[PALU.scala 123:21 136:33]
  wire [63:0] _GEN_157 = io_in_bits_Pctrl_SrcSigned ? _GEN_150 : _GEN_154; // @[PALU.scala 124:28]
  wire [64:0] _T_334 = {_GEN_156,_GEN_157}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_159 = io_in_bits_Pctrl_Translation ? io_in_bits_Pctrl_adderRes_ori[64:1] : io_in_bits_Pctrl_adderRes; // @[PALU.scala 215:32 216:28]
  wire [63:0] _GEN_160 = io_in_bits_Pctrl_Saturating ? _T_334[63:0] : _GEN_159; // @[PALU.scala 211:25 213:28]
  wire  _GEN_161 = io_in_bits_Pctrl_Saturating & _T_334[64]; // @[PALU.scala 211:25 214:21]
  wire [31:0] _T_349 = _T_317[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_350 = {_T_349,_T_317[31:0]}; // @[Cat.scala 30:58]
  wire [80:0] _T_351 = io_in_bits_Pctrl_adderRes_ori + 80'h1; // @[PALU.scala 221:40]
  wire [63:0] _GEN_162 = io_in_bits_Pctrl_isAve ? _T_351[64:1] : io_in_bits_Pctrl_adderRes; // @[PALU.scala 220:22 221:24]
  wire [63:0] _GEN_163 = io_in_bits_Pctrl_isSub_C31 | io_in_bits_Pctrl_isAdd_C31 ? _T_350 : _GEN_162; // @[PALU.scala 218:37 219:24]
  wire [63:0] _GEN_164 = io_in_bits_Pctrl_isAdd_64 | io_in_bits_Pctrl_isSub_64 ? _GEN_160 : _GEN_163; // @[PALU.scala 210:36]
  wire  _GEN_165 = (io_in_bits_Pctrl_isAdd_64 | io_in_bits_Pctrl_isSub_64) & _GEN_161; // @[PALU.scala 210:36]
  wire [63:0] _GEN_166 = io_in_bits_Pctrl_isAdd_32 | io_in_bits_Pctrl_isSub_32 | io_in_bits_Pctrl_isCras_32 |
    io_in_bits_Pctrl_isCrsa_32 | io_in_bits_Pctrl_isStas_32 | io_in_bits_Pctrl_isStsa_32 | io_in_bits_Pctrl_isAdd_Q31 |
    io_in_bits_Pctrl_isSub_Q31 ? _GEN_147 : _GEN_164; // @[PALU.scala 201:108]
  wire  _GEN_167 = io_in_bits_Pctrl_isAdd_32 | io_in_bits_Pctrl_isSub_32 | io_in_bits_Pctrl_isCras_32 |
    io_in_bits_Pctrl_isCrsa_32 | io_in_bits_Pctrl_isStas_32 | io_in_bits_Pctrl_isStsa_32 | io_in_bits_Pctrl_isAdd_Q31 |
    io_in_bits_Pctrl_isSub_Q31 ? _GEN_148 : _GEN_165; // @[PALU.scala 201:108]
  wire [63:0] _GEN_168 = io_in_bits_Pctrl_isAdd_8 | io_in_bits_Pctrl_isSub_8 ? _GEN_124 : _GEN_166; // @[PALU.scala 193:34]
  wire  _GEN_169 = io_in_bits_Pctrl_isAdd_8 | io_in_bits_Pctrl_isSub_8 ? _GEN_125 : _GEN_167; // @[PALU.scala 193:34]
  wire [63:0] adderRes_final = io_in_bits_Pctrl_isAdd_16 | io_in_bits_Pctrl_isSub_16 | io_in_bits_Pctrl_isCras_16 |
    io_in_bits_Pctrl_isCrsa_16 | io_in_bits_Pctrl_isStas_16 | io_in_bits_Pctrl_isStsa_16 | io_in_bits_Pctrl_isAdd_Q15 |
    io_in_bits_Pctrl_isSub_Q15 ? _GEN_41 : _GEN_168; // @[PALU.scala 184:101]
  wire  adderOV = io_in_bits_Pctrl_isAdd_16 | io_in_bits_Pctrl_isSub_16 | io_in_bits_Pctrl_isCras_16 |
    io_in_bits_Pctrl_isCrsa_16 | io_in_bits_Pctrl_isStas_16 | io_in_bits_Pctrl_isStsa_16 | io_in_bits_Pctrl_isAdd_Q15 |
    io_in_bits_Pctrl_isSub_Q15 ? _GEN_42 : _GEN_169; // @[PALU.scala 184:101]
  wire  _T_356 = io_in_bits_Pctrl_adderRes_ori[15:0] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_358 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[16] | _T_356 : _T_356; // @[PALU.scala 164:55]
  wire  _T_359 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[16] : _T_358; // @[PALU.scala 164:31]
  wire [15:0] _T_361 = _T_359 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire  _T_365 = io_in_bits_Pctrl_adderRes_ori[33:18] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_367 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[34] | _T_365 : _T_365; // @[PALU.scala 164:55]
  wire  _T_368 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[34] : _T_367; // @[PALU.scala 164:31]
  wire [15:0] _T_370 = _T_368 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire  _T_374 = io_in_bits_Pctrl_adderRes_ori[51:36] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_376 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[52] | _T_374 : _T_374; // @[PALU.scala 164:55]
  wire  _T_377 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[52] : _T_376; // @[PALU.scala 164:31]
  wire [15:0] _T_379 = _T_377 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire  _T_383 = io_in_bits_Pctrl_adderRes_ori[69:54] == 16'h0; // @[PALU.scala 163:97]
  wire  _T_385 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[70] | _T_383 : _T_383; // @[PALU.scala 164:55]
  wire  _T_386 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[70] : _T_385; // @[PALU.scala 164:31]
  wire [15:0] _T_388 = _T_386 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_391 = {_T_388,_T_379,_T_370,_T_361}; // @[Cat.scala 30:58]
  wire  _T_395 = io_in_bits_Pctrl_adderRes_ori[7:0] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_397 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[8] | _T_395 : _T_395; // @[PALU.scala 164:55]
  wire  _T_398 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[8] : _T_397; // @[PALU.scala 164:31]
  wire [7:0] _T_400 = _T_398 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_404 = io_in_bits_Pctrl_adderRes_ori[17:10] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_406 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[18] | _T_404 : _T_404; // @[PALU.scala 164:55]
  wire  _T_407 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[18] : _T_406; // @[PALU.scala 164:31]
  wire [7:0] _T_409 = _T_407 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_413 = io_in_bits_Pctrl_adderRes_ori[27:20] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_415 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[28] | _T_413 : _T_413; // @[PALU.scala 164:55]
  wire  _T_416 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[28] : _T_415; // @[PALU.scala 164:31]
  wire [7:0] _T_418 = _T_416 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_422 = io_in_bits_Pctrl_adderRes_ori[37:30] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_424 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[38] | _T_422 : _T_422; // @[PALU.scala 164:55]
  wire  _T_425 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[38] : _T_424; // @[PALU.scala 164:31]
  wire [7:0] _T_427 = _T_425 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_431 = io_in_bits_Pctrl_adderRes_ori[47:40] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_433 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[48] | _T_431 : _T_431; // @[PALU.scala 164:55]
  wire  _T_434 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[48] : _T_433; // @[PALU.scala 164:31]
  wire [7:0] _T_436 = _T_434 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_440 = io_in_bits_Pctrl_adderRes_ori[57:50] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_442 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[58] | _T_440 : _T_440; // @[PALU.scala 164:55]
  wire  _T_443 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[58] : _T_442; // @[PALU.scala 164:31]
  wire [7:0] _T_445 = _T_443 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_449 = io_in_bits_Pctrl_adderRes_ori[67:60] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_451 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[68] | _T_449 : _T_449; // @[PALU.scala 164:55]
  wire  _T_452 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[68] : _T_451; // @[PALU.scala 164:31]
  wire [7:0] _T_454 = _T_452 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_458 = io_in_bits_Pctrl_adderRes_ori[77:70] == 8'h0; // @[PALU.scala 163:97]
  wire  _T_460 = io_in_bits_Pctrl_LessEqual ? io_in_bits_Pctrl_adderRes_ori[78] | _T_458 : _T_458; // @[PALU.scala 164:55]
  wire  _T_461 = io_in_bits_Pctrl_LessThan ? io_in_bits_Pctrl_adderRes_ori[78] : _T_460; // @[PALU.scala 164:31]
  wire [7:0] _T_463 = _T_461 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_470 = {_T_463,_T_454,_T_445,_T_436,_T_427,_T_418,_T_409,_T_400}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_172 = io_in_bits_Pctrl_isComp_8 ? _T_470 : 64'h0; // @[PALU.scala 228:25 229:20]
  wire [63:0] compareRes = io_in_bits_Pctrl_isComp_16 ? _T_391 : _GEN_172; // @[PALU.scala 226:20 227:20]
  wire  _T_473 = ~io_in_bits_DecodeIn_ctrl_fuOpType[0]; // @[PALU.scala 235:55]
  wire [15:0] _T_480 = ~(io_in_bits_Pctrl_adderRes_ori[16] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[15:0] :
    io_in_bits_DecodeIn_data_src2[15:0]; // @[PALU.scala 175:30]
  wire [15:0] _T_498 = ~(io_in_bits_Pctrl_adderRes_ori[34] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[31:16] :
    io_in_bits_DecodeIn_data_src2[31:16]; // @[PALU.scala 175:30]
  wire [15:0] _T_516 = ~(io_in_bits_Pctrl_adderRes_ori[52] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[47:32] :
    io_in_bits_DecodeIn_data_src2[47:32]; // @[PALU.scala 175:30]
  wire [15:0] _T_534 = ~(io_in_bits_Pctrl_adderRes_ori[70] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[63:48] :
    io_in_bits_DecodeIn_data_src2[63:48]; // @[PALU.scala 175:30]
  wire [63:0] _T_548 = {_T_534,_T_516,_T_498,_T_480}; // @[Cat.scala 30:58]
  wire [7:0] _T_558 = ~(io_in_bits_Pctrl_adderRes_ori[8] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src2[7:0]; // @[PALU.scala 175:30]
  wire [7:0] _T_576 = ~(io_in_bits_Pctrl_adderRes_ori[18] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[15:8] :
    io_in_bits_DecodeIn_data_src2[15:8]; // @[PALU.scala 175:30]
  wire [7:0] _T_594 = ~(io_in_bits_Pctrl_adderRes_ori[28] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[23:16] :
    io_in_bits_DecodeIn_data_src2[23:16]; // @[PALU.scala 175:30]
  wire [7:0] _T_612 = ~(io_in_bits_Pctrl_adderRes_ori[38] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[31:24] :
    io_in_bits_DecodeIn_data_src2[31:24]; // @[PALU.scala 175:30]
  wire [7:0] _T_630 = ~(io_in_bits_Pctrl_adderRes_ori[48] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[39:32] :
    io_in_bits_DecodeIn_data_src2[39:32]; // @[PALU.scala 175:30]
  wire [7:0] _T_648 = ~(io_in_bits_Pctrl_adderRes_ori[58] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[47:40] :
    io_in_bits_DecodeIn_data_src2[47:40]; // @[PALU.scala 175:30]
  wire [7:0] _T_666 = ~(io_in_bits_Pctrl_adderRes_ori[68] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[55:48] :
    io_in_bits_DecodeIn_data_src2[55:48]; // @[PALU.scala 175:30]
  wire [7:0] _T_684 = ~(io_in_bits_Pctrl_adderRes_ori[78] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[63:56] :
    io_in_bits_DecodeIn_data_src2[63:56]; // @[PALU.scala 175:30]
  wire [63:0] _T_702 = {_T_684,_T_666,_T_648,_T_630,_T_612,_T_594,_T_576,_T_558}; // @[Cat.scala 30:58]
  wire  _T_705 = ~io_in_bits_DecodeIn_ctrl_funct3[1]; // @[PALU.scala 239:58]
  wire [63:0] _T_712 = ~(io_in_bits_Pctrl_adderRes_ori[64] ^ _T_705) ? io_in_bits_DecodeIn_data_src1 :
    io_in_bits_DecodeIn_data_src2; // @[PALU.scala 175:30]
  wire [31:0] _T_733 = ~(io_in_bits_Pctrl_adderRes_ori[32] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[31:0] :
    io_in_bits_DecodeIn_data_src2[31:0]; // @[PALU.scala 175:30]
  wire [31:0] _T_751 = ~(io_in_bits_Pctrl_adderRes_ori[66] ^ _T_473) ? io_in_bits_DecodeIn_data_src1[63:32] :
    io_in_bits_DecodeIn_data_src2[63:32]; // @[PALU.scala 175:30]
  wire [63:0] _T_763 = {_T_751,_T_733}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_174 = io_in_bits_Pctrl_isMaxMin_32 ? _T_763 : 64'h0; // @[PALU.scala 240:28 241:19]
  wire [63:0] _GEN_175 = io_in_bits_Pctrl_isMaxMin_XLEN ? _T_712 : _GEN_174; // @[PALU.scala 238:30 239:19]
  wire [63:0] _GEN_176 = io_in_bits_Pctrl_isMaxMin_8 ? _T_702 : _GEN_175; // @[PALU.scala 236:27 237:19]
  wire [63:0] maxminRes = io_in_bits_Pctrl_isMaxMin_16 ? _T_548 : _GEN_176; // @[PALU.scala 234:22 235:19]
  wire [63:0] _T_766 = io_in_bits_DecodeIn_ctrl_fuOpType[0] ? io_in_bits_DecodeIn_data_src3 : 64'h0; // @[PALU.scala 247:22]
  wire [7:0] _T_770 = 8'hff ^ io_in_bits_Pctrl_adderRes[7:0]; // @[PALU.scala 247:128]
  wire [7:0] _T_772 = _T_770 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_774 = io_in_bits_Pctrl_adderRes_ori[8] ? _T_772 : io_in_bits_Pctrl_adderRes[7:0]; // @[PALU.scala 247:79]
  wire [7:0] _T_778 = 8'hff ^ io_in_bits_Pctrl_adderRes[15:8]; // @[PALU.scala 247:128]
  wire [7:0] _T_780 = _T_778 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_782 = io_in_bits_Pctrl_adderRes_ori[18] ? _T_780 : io_in_bits_Pctrl_adderRes[15:8]; // @[PALU.scala 247:79]
  wire [7:0] _T_786 = 8'hff ^ io_in_bits_Pctrl_adderRes[23:16]; // @[PALU.scala 247:128]
  wire [7:0] _T_788 = _T_786 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_790 = io_in_bits_Pctrl_adderRes_ori[28] ? _T_788 : io_in_bits_Pctrl_adderRes[23:16]; // @[PALU.scala 247:79]
  wire [7:0] _T_794 = 8'hff ^ io_in_bits_Pctrl_adderRes[31:24]; // @[PALU.scala 247:128]
  wire [7:0] _T_796 = _T_794 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_798 = io_in_bits_Pctrl_adderRes_ori[38] ? _T_796 : io_in_bits_Pctrl_adderRes[31:24]; // @[PALU.scala 247:79]
  wire [7:0] _T_802 = 8'hff ^ io_in_bits_Pctrl_adderRes[39:32]; // @[PALU.scala 247:128]
  wire [7:0] _T_804 = _T_802 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_806 = io_in_bits_Pctrl_adderRes_ori[48] ? _T_804 : io_in_bits_Pctrl_adderRes[39:32]; // @[PALU.scala 247:79]
  wire [7:0] _T_810 = 8'hff ^ io_in_bits_Pctrl_adderRes[47:40]; // @[PALU.scala 247:128]
  wire [7:0] _T_812 = _T_810 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_814 = io_in_bits_Pctrl_adderRes_ori[58] ? _T_812 : io_in_bits_Pctrl_adderRes[47:40]; // @[PALU.scala 247:79]
  wire [7:0] _T_818 = 8'hff ^ io_in_bits_Pctrl_adderRes[55:48]; // @[PALU.scala 247:128]
  wire [7:0] _T_820 = _T_818 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_822 = io_in_bits_Pctrl_adderRes_ori[68] ? _T_820 : io_in_bits_Pctrl_adderRes[55:48]; // @[PALU.scala 247:79]
  wire [7:0] _T_826 = 8'hff ^ io_in_bits_Pctrl_adderRes[63:56]; // @[PALU.scala 247:128]
  wire [7:0] _T_828 = _T_826 + 8'h1; // @[PALU.scala 247:151]
  wire [7:0] _T_830 = io_in_bits_Pctrl_adderRes_ori[78] ? _T_828 : io_in_bits_Pctrl_adderRes[63:56]; // @[PALU.scala 247:79]
  wire [8:0] _T_831 = _T_774 + _T_782; // @[PALU.scala 247:188]
  wire [8:0] _GEN_648 = {{1'd0}, _T_790}; // @[PALU.scala 247:188]
  wire [9:0] _T_832 = _T_831 + _GEN_648; // @[PALU.scala 247:188]
  wire [9:0] _GEN_649 = {{2'd0}, _T_798}; // @[PALU.scala 247:188]
  wire [10:0] _T_833 = _T_832 + _GEN_649; // @[PALU.scala 247:188]
  wire [10:0] _GEN_650 = {{3'd0}, _T_806}; // @[PALU.scala 247:188]
  wire [11:0] _T_834 = _T_833 + _GEN_650; // @[PALU.scala 247:188]
  wire [11:0] _GEN_651 = {{4'd0}, _T_814}; // @[PALU.scala 247:188]
  wire [12:0] _T_835 = _T_834 + _GEN_651; // @[PALU.scala 247:188]
  wire [12:0] _GEN_652 = {{5'd0}, _T_822}; // @[PALU.scala 247:188]
  wire [13:0] _T_836 = _T_835 + _GEN_652; // @[PALU.scala 247:188]
  wire [13:0] _GEN_653 = {{6'd0}, _T_830}; // @[PALU.scala 247:188]
  wire [14:0] _T_837 = _T_836 + _GEN_653; // @[PALU.scala 247:188]
  wire [63:0] _GEN_654 = {{49'd0}, _T_837}; // @[PALU.scala 247:48]
  wire [63:0] _T_839 = _T_766 + _GEN_654; // @[PALU.scala 247:48]
  wire [63:0] pbsRes = io_in_bits_Pctrl_isPbs ? _T_839 : 64'h0; // @[PALU.scala 246:16 247:16]
  wire [4:0] _T_875 = 5'h1f ^ io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 367:52]
  wire [4:0] _T_877 = _T_875 + 5'h1; // @[PALU.scala 367:79]
  wire [4:0] _GEN_179 = _T_877 == 5'h10 ? 5'hf : _T_877; // @[PALU.scala 368:26 369:65 370:30]
  wire [4:0] _GEN_180 = io_in_bits_DecodeIn_data_src2[4] ? _GEN_179 : io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 366:47]
  wire [5:0] _T_884 = {io_in_bits_DecodeIn_data_src2[4],_GEN_180}; // @[Cat.scala 30:58]
  wire [3:0] _T_890 = 4'hf ^ io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 367:52]
  wire [3:0] _T_892 = _T_890 + 4'h1; // @[PALU.scala 367:79]
  wire [3:0] _GEN_182 = _T_892 == 4'h8 ? 4'h7 : _T_892; // @[PALU.scala 368:26 369:65 370:30]
  wire [3:0] _GEN_183 = io_in_bits_DecodeIn_data_src2[3] ? _GEN_182 : io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 366:47]
  wire [4:0] _T_899 = {io_in_bits_DecodeIn_data_src2[3],io_in_bits_DecodeIn_data_src2[3:0]}; // @[Cat.scala 30:58]
  wire [5:0] _T_900 = io_in_bits_Pctrl_isLR_16 ? _T_884 : {{1'd0}, _T_899}; // @[PALU.scala 500:22]
  wire [63:0] _WIRE_80 = {{58'd0}, _T_900};
  wire [4:0] _T_903 = io_in_bits_Pctrl_isLR_16 ? _WIRE_80[4:0] : {{1'd0}, _WIRE_80[3:0]}; // @[PALU.scala 501:27]
  wire  _T_907 = io_in_bits_Pctrl_isRs_16 | io_in_bits_Pctrl_isLR_16 & _WIRE_80[5]; // @[PALU.scala 503:70]
  wire [4:0] _T_911 = _T_903 - 5'h1; // @[PALU.scala 327:50]
  wire [4:0] _GEN_185 = io_in_bits_Pctrl_Round ? _T_911 : _T_903; // @[PALU.scala 327:{32,42}]
  wire [15:0] _T_912 = io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 329:42]
  wire [15:0] _T_914 = $signed(_T_912) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_915 = io_in_bits_DecodeIn_data_src1[15:0] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_186 = io_in_bits_Pctrl_Arithmetic ? _T_914 : _T_915; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_917 = {_GEN_186[15],_GEN_186}; // @[Cat.scala 30:58]
  wire [16:0] _T_918 = {1'h0,_GEN_186}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_187 = io_in_bits_Pctrl_Arithmetic ? _T_917 : _T_918; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_920 = _GEN_187 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_188 = io_in_bits_Pctrl_Round ? _T_920[16:1] : _GEN_186; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_931 = io_in_bits_DecodeIn_data_src1[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_932 = {_T_931,io_in_bits_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_2 = {{31'd0}, _T_932}; // @[PALU.scala 341:35]
  wire [62:0] _T_933 = _GEN_2 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_938 = 63'hffffffff ^ _T_933; // @[PALU.scala 345:80]
  wire [62:0] _GEN_189 = _T_933[31] ? _T_938 : _T_933; // @[PALU.scala 345:{53,59}]
  wire  _T_940 = _GEN_189[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_190 = _T_933[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_192 = _GEN_189[31:15] != 17'h0 ? _GEN_190 : _T_933[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_193 = io_in_bits_Pctrl_ShiftSigned & _T_940; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_194 = io_in_bits_Pctrl_ShiftSigned ? _GEN_192 : _T_933[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_195 = _T_907 ? _GEN_188 : _GEN_194; // @[PALU.scala 323:32]
  wire  _GEN_196 = _T_907 ? 1'h0 : _GEN_193; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_197 = _T_903 != 5'h0 ? _GEN_195 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_198 = _T_903 != 5'h0 & _GEN_196; // @[PALU.scala 322:31 317:45]
  wire [15:0] _T_966 = io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 329:42]
  wire [15:0] _T_968 = $signed(_T_966) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_969 = io_in_bits_DecodeIn_data_src1[31:16] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_200 = io_in_bits_Pctrl_Arithmetic ? _T_968 : _T_969; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_971 = {_GEN_200[15],_GEN_200}; // @[Cat.scala 30:58]
  wire [16:0] _T_972 = {1'h0,_GEN_200}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_201 = io_in_bits_Pctrl_Arithmetic ? _T_971 : _T_972; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_974 = _GEN_201 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_202 = io_in_bits_Pctrl_Round ? _T_974[16:1] : _GEN_200; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_985 = io_in_bits_DecodeIn_data_src1[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_986 = {_T_985,io_in_bits_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_4 = {{31'd0}, _T_986}; // @[PALU.scala 341:35]
  wire [62:0] _T_987 = _GEN_4 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_992 = 63'hffffffff ^ _T_987; // @[PALU.scala 345:80]
  wire [62:0] _GEN_203 = _T_987[31] ? _T_992 : _T_987; // @[PALU.scala 345:{53,59}]
  wire  _T_994 = _GEN_203[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_204 = _T_987[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_206 = _GEN_203[31:15] != 17'h0 ? _GEN_204 : _T_987[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_207 = io_in_bits_Pctrl_ShiftSigned & _T_994; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_208 = io_in_bits_Pctrl_ShiftSigned ? _GEN_206 : _T_987[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_209 = _T_907 ? _GEN_202 : _GEN_208; // @[PALU.scala 323:32]
  wire  _GEN_210 = _T_907 ? 1'h0 : _GEN_207; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_211 = _T_903 != 5'h0 ? _GEN_209 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_212 = _T_903 != 5'h0 & _GEN_210; // @[PALU.scala 322:31 317:45]
  wire [15:0] _T_1020 = io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 329:42]
  wire [15:0] _T_1022 = $signed(_T_1020) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_1023 = io_in_bits_DecodeIn_data_src1[47:32] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_214 = io_in_bits_Pctrl_Arithmetic ? _T_1022 : _T_1023; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_1025 = {_GEN_214[15],_GEN_214}; // @[Cat.scala 30:58]
  wire [16:0] _T_1026 = {1'h0,_GEN_214}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_215 = io_in_bits_Pctrl_Arithmetic ? _T_1025 : _T_1026; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_1028 = _GEN_215 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_216 = io_in_bits_Pctrl_Round ? _T_1028[16:1] : _GEN_214; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_1039 = io_in_bits_DecodeIn_data_src1[47] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1040 = {_T_1039,io_in_bits_DecodeIn_data_src1[47:32]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_6 = {{31'd0}, _T_1040}; // @[PALU.scala 341:35]
  wire [62:0] _T_1041 = _GEN_6 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_1046 = 63'hffffffff ^ _T_1041; // @[PALU.scala 345:80]
  wire [62:0] _GEN_217 = _T_1041[31] ? _T_1046 : _T_1041; // @[PALU.scala 345:{53,59}]
  wire  _T_1048 = _GEN_217[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_218 = _T_1041[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_220 = _GEN_217[31:15] != 17'h0 ? _GEN_218 : _T_1041[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_221 = io_in_bits_Pctrl_ShiftSigned & _T_1048; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_222 = io_in_bits_Pctrl_ShiftSigned ? _GEN_220 : _T_1041[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_223 = _T_907 ? _GEN_216 : _GEN_222; // @[PALU.scala 323:32]
  wire  _GEN_224 = _T_907 ? 1'h0 : _GEN_221; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_225 = _T_903 != 5'h0 ? _GEN_223 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_226 = _T_903 != 5'h0 & _GEN_224; // @[PALU.scala 322:31 317:45]
  wire [15:0] _T_1074 = io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 329:42]
  wire [15:0] _T_1076 = $signed(_T_1074) >>> _GEN_185; // @[PALU.scala 329:62]
  wire [15:0] _T_1077 = io_in_bits_DecodeIn_data_src1[63:48] >> _GEN_185; // @[PALU.scala 331:41]
  wire [15:0] _GEN_228 = io_in_bits_Pctrl_Arithmetic ? _T_1076 : _T_1077; // @[PALU.scala 328:37 329:29 331:29]
  wire [16:0] _T_1079 = {_GEN_228[15],_GEN_228}; // @[Cat.scala 30:58]
  wire [16:0] _T_1080 = {1'h0,_GEN_228}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_229 = io_in_bits_Pctrl_Arithmetic ? _T_1079 : _T_1080; // @[PALU.scala 96:24 97:15 99:15]
  wire [16:0] _T_1082 = _GEN_229 + 17'h1; // @[PALU.scala 334:66]
  wire [15:0] _GEN_230 = io_in_bits_Pctrl_Round ? _T_1082[16:1] : _GEN_228; // @[PALU.scala 333:32 334:29 336:29]
  wire [15:0] _T_1093 = io_in_bits_DecodeIn_data_src1[63] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1094 = {_T_1093,io_in_bits_DecodeIn_data_src1[63:48]}; // @[Cat.scala 30:58]
  wire [62:0] _GEN_9 = {{31'd0}, _T_1094}; // @[PALU.scala 341:35]
  wire [62:0] _T_1095 = _GEN_9 << _T_903; // @[PALU.scala 341:35]
  wire [62:0] _T_1100 = 63'hffffffff ^ _T_1095; // @[PALU.scala 345:80]
  wire [62:0] _GEN_231 = _T_1095[31] ? _T_1100 : _T_1095; // @[PALU.scala 345:{53,59}]
  wire  _T_1102 = _GEN_231[31:15] != 17'h0; // @[PALU.scala 346:54]
  wire [15:0] _GEN_232 = _T_1095[31] ? 16'h8000 : 16'h7fff; // @[PALU.scala 348:57 349:37 351:37]
  wire [15:0] _GEN_234 = _GEN_231[31:15] != 17'h0 ? _GEN_232 : _T_1095[15:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_235 = io_in_bits_Pctrl_ShiftSigned & _T_1102; // @[PALU.scala 343:38 317:45]
  wire [15:0] _GEN_236 = io_in_bits_Pctrl_ShiftSigned ? _GEN_234 : _T_1095[15:0]; // @[PALU.scala 342:25 343:38]
  wire [15:0] _GEN_237 = _T_907 ? _GEN_230 : _GEN_236; // @[PALU.scala 323:32]
  wire  _GEN_238 = _T_907 ? 1'h0 : _GEN_235; // @[PALU.scala 323:32 317:45]
  wire [15:0] _GEN_239 = _T_903 != 5'h0 ? _GEN_237 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_240 = _T_903 != 5'h0 & _GEN_238; // @[PALU.scala 322:31 317:45]
  wire  _T_1126 = _GEN_198 | _GEN_212 | _GEN_226 | _GEN_240; // @[PALU.scala 361:24]
  wire [64:0] _T_1130 = {_T_1126,_GEN_239,_GEN_225,_GEN_211,_GEN_197}; // @[Cat.scala 30:58]
  wire [4:0] _T_1150 = {io_in_bits_DecodeIn_data_src2[3],_GEN_183}; // @[Cat.scala 30:58]
  wire [3:0] _T_1165 = {io_in_bits_DecodeIn_data_src2[2],io_in_bits_DecodeIn_data_src2[2:0]}; // @[Cat.scala 30:58]
  wire [4:0] _T_1166 = io_in_bits_Pctrl_isLR_8 ? _T_1150 : {{1'd0}, _T_1165}; // @[PALU.scala 508:22]
  wire [63:0] _WIRE_120 = {{59'd0}, _T_1166};
  wire [3:0] _T_1169 = io_in_bits_Pctrl_isLR_8 ? _WIRE_120[3:0] : {{1'd0}, _WIRE_120[2:0]}; // @[PALU.scala 509:27]
  wire  _T_1173 = io_in_bits_Pctrl_isRs_8 | io_in_bits_Pctrl_isLR_8 & _WIRE_120[4]; // @[PALU.scala 511:68]
  wire [3:0] _T_1177 = _T_1169 - 4'h1; // @[PALU.scala 327:50]
  wire [3:0] _GEN_247 = io_in_bits_Pctrl_Round ? _T_1177 : _T_1169; // @[PALU.scala 327:{32,42}]
  wire [7:0] _T_1178 = io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 329:42]
  wire [7:0] _T_1180 = $signed(_T_1178) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1181 = io_in_bits_DecodeIn_data_src1[7:0] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_248 = io_in_bits_Pctrl_Arithmetic ? _T_1180 : _T_1181; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1183 = {_GEN_248[7],_GEN_248}; // @[Cat.scala 30:58]
  wire [8:0] _T_1184 = {1'h0,_GEN_248}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_249 = io_in_bits_Pctrl_Arithmetic ? _T_1183 : _T_1184; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1186 = _GEN_249 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_250 = io_in_bits_Pctrl_Round ? _T_1186[8:1] : _GEN_248; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1197 = io_in_bits_DecodeIn_data_src1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1198 = {_T_1197,io_in_bits_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_14 = {{15'd0}, _T_1198}; // @[PALU.scala 341:35]
  wire [30:0] _T_1199 = _GEN_14 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1204 = 31'hffff ^ _T_1199; // @[PALU.scala 345:80]
  wire [30:0] _GEN_251 = _T_1199[15] ? _T_1204 : _T_1199; // @[PALU.scala 345:{53,59}]
  wire  _T_1206 = _GEN_251[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_252 = _T_1199[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_254 = _GEN_251[15:7] != 9'h0 ? _GEN_252 : _T_1199[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_255 = io_in_bits_Pctrl_ShiftSigned & _T_1206; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_256 = io_in_bits_Pctrl_ShiftSigned ? _GEN_254 : _T_1199[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_257 = _T_1173 ? _GEN_250 : _GEN_256; // @[PALU.scala 323:32]
  wire  _GEN_258 = _T_1173 ? 1'h0 : _GEN_255; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_259 = _T_1169 != 4'h0 ? _GEN_257 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_260 = _T_1169 != 4'h0 & _GEN_258; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1232 = io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 329:42]
  wire [7:0] _T_1234 = $signed(_T_1232) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1235 = io_in_bits_DecodeIn_data_src1[15:8] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_262 = io_in_bits_Pctrl_Arithmetic ? _T_1234 : _T_1235; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1237 = {_GEN_262[7],_GEN_262}; // @[Cat.scala 30:58]
  wire [8:0] _T_1238 = {1'h0,_GEN_262}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_263 = io_in_bits_Pctrl_Arithmetic ? _T_1237 : _T_1238; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1240 = _GEN_263 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_264 = io_in_bits_Pctrl_Round ? _T_1240[8:1] : _GEN_262; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1251 = io_in_bits_DecodeIn_data_src1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1252 = {_T_1251,io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_16 = {{15'd0}, _T_1252}; // @[PALU.scala 341:35]
  wire [30:0] _T_1253 = _GEN_16 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1258 = 31'hffff ^ _T_1253; // @[PALU.scala 345:80]
  wire [30:0] _GEN_265 = _T_1253[15] ? _T_1258 : _T_1253; // @[PALU.scala 345:{53,59}]
  wire  _T_1260 = _GEN_265[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_266 = _T_1253[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_268 = _GEN_265[15:7] != 9'h0 ? _GEN_266 : _T_1253[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_269 = io_in_bits_Pctrl_ShiftSigned & _T_1260; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_270 = io_in_bits_Pctrl_ShiftSigned ? _GEN_268 : _T_1253[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_271 = _T_1173 ? _GEN_264 : _GEN_270; // @[PALU.scala 323:32]
  wire  _GEN_272 = _T_1173 ? 1'h0 : _GEN_269; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_273 = _T_1169 != 4'h0 ? _GEN_271 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_274 = _T_1169 != 4'h0 & _GEN_272; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1286 = io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 329:42]
  wire [7:0] _T_1288 = $signed(_T_1286) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1289 = io_in_bits_DecodeIn_data_src1[23:16] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_276 = io_in_bits_Pctrl_Arithmetic ? _T_1288 : _T_1289; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1291 = {_GEN_276[7],_GEN_276}; // @[Cat.scala 30:58]
  wire [8:0] _T_1292 = {1'h0,_GEN_276}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_277 = io_in_bits_Pctrl_Arithmetic ? _T_1291 : _T_1292; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1294 = _GEN_277 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_278 = io_in_bits_Pctrl_Round ? _T_1294[8:1] : _GEN_276; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1305 = io_in_bits_DecodeIn_data_src1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1306 = {_T_1305,io_in_bits_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_24 = {{15'd0}, _T_1306}; // @[PALU.scala 341:35]
  wire [30:0] _T_1307 = _GEN_24 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1312 = 31'hffff ^ _T_1307; // @[PALU.scala 345:80]
  wire [30:0] _GEN_279 = _T_1307[15] ? _T_1312 : _T_1307; // @[PALU.scala 345:{53,59}]
  wire  _T_1314 = _GEN_279[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_280 = _T_1307[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_282 = _GEN_279[15:7] != 9'h0 ? _GEN_280 : _T_1307[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_283 = io_in_bits_Pctrl_ShiftSigned & _T_1314; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_284 = io_in_bits_Pctrl_ShiftSigned ? _GEN_282 : _T_1307[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_285 = _T_1173 ? _GEN_278 : _GEN_284; // @[PALU.scala 323:32]
  wire  _GEN_286 = _T_1173 ? 1'h0 : _GEN_283; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_287 = _T_1169 != 4'h0 ? _GEN_285 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_288 = _T_1169 != 4'h0 & _GEN_286; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1340 = io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 329:42]
  wire [7:0] _T_1342 = $signed(_T_1340) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1343 = io_in_bits_DecodeIn_data_src1[31:24] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_290 = io_in_bits_Pctrl_Arithmetic ? _T_1342 : _T_1343; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1345 = {_GEN_290[7],_GEN_290}; // @[Cat.scala 30:58]
  wire [8:0] _T_1346 = {1'h0,_GEN_290}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_291 = io_in_bits_Pctrl_Arithmetic ? _T_1345 : _T_1346; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1348 = _GEN_291 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_292 = io_in_bits_Pctrl_Round ? _T_1348[8:1] : _GEN_290; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1359 = io_in_bits_DecodeIn_data_src1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1360 = {_T_1359,io_in_bits_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_26 = {{15'd0}, _T_1360}; // @[PALU.scala 341:35]
  wire [30:0] _T_1361 = _GEN_26 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1366 = 31'hffff ^ _T_1361; // @[PALU.scala 345:80]
  wire [30:0] _GEN_293 = _T_1361[15] ? _T_1366 : _T_1361; // @[PALU.scala 345:{53,59}]
  wire  _T_1368 = _GEN_293[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_294 = _T_1361[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_296 = _GEN_293[15:7] != 9'h0 ? _GEN_294 : _T_1361[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_297 = io_in_bits_Pctrl_ShiftSigned & _T_1368; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_298 = io_in_bits_Pctrl_ShiftSigned ? _GEN_296 : _T_1361[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_299 = _T_1173 ? _GEN_292 : _GEN_298; // @[PALU.scala 323:32]
  wire  _GEN_300 = _T_1173 ? 1'h0 : _GEN_297; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_301 = _T_1169 != 4'h0 ? _GEN_299 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_302 = _T_1169 != 4'h0 & _GEN_300; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1394 = io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 329:42]
  wire [7:0] _T_1396 = $signed(_T_1394) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1397 = io_in_bits_DecodeIn_data_src1[39:32] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_304 = io_in_bits_Pctrl_Arithmetic ? _T_1396 : _T_1397; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1399 = {_GEN_304[7],_GEN_304}; // @[Cat.scala 30:58]
  wire [8:0] _T_1400 = {1'h0,_GEN_304}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_305 = io_in_bits_Pctrl_Arithmetic ? _T_1399 : _T_1400; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1402 = _GEN_305 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_306 = io_in_bits_Pctrl_Round ? _T_1402[8:1] : _GEN_304; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1413 = io_in_bits_DecodeIn_data_src1[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1414 = {_T_1413,io_in_bits_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_34 = {{15'd0}, _T_1414}; // @[PALU.scala 341:35]
  wire [30:0] _T_1415 = _GEN_34 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1420 = 31'hffff ^ _T_1415; // @[PALU.scala 345:80]
  wire [30:0] _GEN_307 = _T_1415[15] ? _T_1420 : _T_1415; // @[PALU.scala 345:{53,59}]
  wire  _T_1422 = _GEN_307[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_308 = _T_1415[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_310 = _GEN_307[15:7] != 9'h0 ? _GEN_308 : _T_1415[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_311 = io_in_bits_Pctrl_ShiftSigned & _T_1422; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_312 = io_in_bits_Pctrl_ShiftSigned ? _GEN_310 : _T_1415[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_313 = _T_1173 ? _GEN_306 : _GEN_312; // @[PALU.scala 323:32]
  wire  _GEN_314 = _T_1173 ? 1'h0 : _GEN_311; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_315 = _T_1169 != 4'h0 ? _GEN_313 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_316 = _T_1169 != 4'h0 & _GEN_314; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1448 = io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 329:42]
  wire [7:0] _T_1450 = $signed(_T_1448) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1451 = io_in_bits_DecodeIn_data_src1[47:40] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_318 = io_in_bits_Pctrl_Arithmetic ? _T_1450 : _T_1451; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1453 = {_GEN_318[7],_GEN_318}; // @[Cat.scala 30:58]
  wire [8:0] _T_1454 = {1'h0,_GEN_318}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_319 = io_in_bits_Pctrl_Arithmetic ? _T_1453 : _T_1454; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1456 = _GEN_319 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_320 = io_in_bits_Pctrl_Round ? _T_1456[8:1] : _GEN_318; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1467 = io_in_bits_DecodeIn_data_src1[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1468 = {_T_1467,io_in_bits_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_36 = {{15'd0}, _T_1468}; // @[PALU.scala 341:35]
  wire [30:0] _T_1469 = _GEN_36 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1474 = 31'hffff ^ _T_1469; // @[PALU.scala 345:80]
  wire [30:0] _GEN_321 = _T_1469[15] ? _T_1474 : _T_1469; // @[PALU.scala 345:{53,59}]
  wire  _T_1476 = _GEN_321[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_322 = _T_1469[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_324 = _GEN_321[15:7] != 9'h0 ? _GEN_322 : _T_1469[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_325 = io_in_bits_Pctrl_ShiftSigned & _T_1476; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_326 = io_in_bits_Pctrl_ShiftSigned ? _GEN_324 : _T_1469[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_327 = _T_1173 ? _GEN_320 : _GEN_326; // @[PALU.scala 323:32]
  wire  _GEN_328 = _T_1173 ? 1'h0 : _GEN_325; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_329 = _T_1169 != 4'h0 ? _GEN_327 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_330 = _T_1169 != 4'h0 & _GEN_328; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1502 = io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 329:42]
  wire [7:0] _T_1504 = $signed(_T_1502) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1505 = io_in_bits_DecodeIn_data_src1[55:48] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_332 = io_in_bits_Pctrl_Arithmetic ? _T_1504 : _T_1505; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1507 = {_GEN_332[7],_GEN_332}; // @[Cat.scala 30:58]
  wire [8:0] _T_1508 = {1'h0,_GEN_332}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_333 = io_in_bits_Pctrl_Arithmetic ? _T_1507 : _T_1508; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1510 = _GEN_333 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_334 = io_in_bits_Pctrl_Round ? _T_1510[8:1] : _GEN_332; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1521 = io_in_bits_DecodeIn_data_src1[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1522 = {_T_1521,io_in_bits_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_45 = {{15'd0}, _T_1522}; // @[PALU.scala 341:35]
  wire [30:0] _T_1523 = _GEN_45 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1528 = 31'hffff ^ _T_1523; // @[PALU.scala 345:80]
  wire [30:0] _GEN_335 = _T_1523[15] ? _T_1528 : _T_1523; // @[PALU.scala 345:{53,59}]
  wire  _T_1530 = _GEN_335[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_336 = _T_1523[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_338 = _GEN_335[15:7] != 9'h0 ? _GEN_336 : _T_1523[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_339 = io_in_bits_Pctrl_ShiftSigned & _T_1530; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_340 = io_in_bits_Pctrl_ShiftSigned ? _GEN_338 : _T_1523[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_341 = _T_1173 ? _GEN_334 : _GEN_340; // @[PALU.scala 323:32]
  wire  _GEN_342 = _T_1173 ? 1'h0 : _GEN_339; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_343 = _T_1169 != 4'h0 ? _GEN_341 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_344 = _T_1169 != 4'h0 & _GEN_342; // @[PALU.scala 322:31 317:45]
  wire [7:0] _T_1556 = io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 329:42]
  wire [7:0] _T_1558 = $signed(_T_1556) >>> _GEN_247; // @[PALU.scala 329:62]
  wire [7:0] _T_1559 = io_in_bits_DecodeIn_data_src1[63:56] >> _GEN_247; // @[PALU.scala 331:41]
  wire [7:0] _GEN_346 = io_in_bits_Pctrl_Arithmetic ? _T_1558 : _T_1559; // @[PALU.scala 328:37 329:29 331:29]
  wire [8:0] _T_1561 = {_GEN_346[7],_GEN_346}; // @[Cat.scala 30:58]
  wire [8:0] _T_1562 = {1'h0,_GEN_346}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_347 = io_in_bits_Pctrl_Arithmetic ? _T_1561 : _T_1562; // @[PALU.scala 96:24 97:15 99:15]
  wire [8:0] _T_1564 = _GEN_347 + 9'h1; // @[PALU.scala 334:66]
  wire [7:0] _GEN_348 = io_in_bits_Pctrl_Round ? _T_1564[8:1] : _GEN_346; // @[PALU.scala 333:32 334:29 336:29]
  wire [7:0] _T_1575 = io_in_bits_DecodeIn_data_src1[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1576 = {_T_1575,io_in_bits_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_47 = {{15'd0}, _T_1576}; // @[PALU.scala 341:35]
  wire [30:0] _T_1577 = _GEN_47 << _T_1169; // @[PALU.scala 341:35]
  wire [30:0] _T_1582 = 31'hffff ^ _T_1577; // @[PALU.scala 345:80]
  wire [30:0] _GEN_349 = _T_1577[15] ? _T_1582 : _T_1577; // @[PALU.scala 345:{53,59}]
  wire  _T_1584 = _GEN_349[15:7] != 9'h0; // @[PALU.scala 346:54]
  wire [7:0] _GEN_350 = _T_1577[15] ? 8'h80 : 8'h7f; // @[PALU.scala 348:57 349:37 351:37]
  wire [7:0] _GEN_352 = _GEN_349[15:7] != 9'h0 ? _GEN_350 : _T_1577[7:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_353 = io_in_bits_Pctrl_ShiftSigned & _T_1584; // @[PALU.scala 343:38 317:45]
  wire [7:0] _GEN_354 = io_in_bits_Pctrl_ShiftSigned ? _GEN_352 : _T_1577[7:0]; // @[PALU.scala 342:25 343:38]
  wire [7:0] _GEN_355 = _T_1173 ? _GEN_348 : _GEN_354; // @[PALU.scala 323:32]
  wire  _GEN_356 = _T_1173 ? 1'h0 : _GEN_353; // @[PALU.scala 323:32 317:45]
  wire [7:0] _GEN_357 = _T_1169 != 4'h0 ? _GEN_355 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_358 = _T_1169 != 4'h0 & _GEN_356; // @[PALU.scala 322:31 317:45]
  wire  _T_1612 = _GEN_260 | _GEN_274 | _GEN_288 | _GEN_302 | _GEN_316 | _GEN_330 | _GEN_344 | _GEN_358; // @[PALU.scala 361:24]
  wire [64:0] _T_1620 = {_T_1612,_GEN_357,_GEN_343,_GEN_329,_GEN_315,_GEN_301,_GEN_287,_GEN_273,_GEN_259}; // @[Cat.scala 30:58]
  wire  _T_1636 = io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isLR_32; // @[PALU.scala 517:32]
  wire [5:0] _T_1642 = 6'h3f ^ io_in_bits_DecodeIn_data_src2[5:0]; // @[PALU.scala 367:52]
  wire [5:0] _T_1644 = _T_1642 + 6'h1; // @[PALU.scala 367:79]
  wire [5:0] _GEN_359 = _T_1644 == 6'h20 ? 6'h1f : _T_1644; // @[PALU.scala 368:26 369:65 370:30]
  wire [5:0] _GEN_360 = io_in_bits_DecodeIn_data_src2[5] ? _GEN_359 : io_in_bits_DecodeIn_data_src2[5:0]; // @[PALU.scala 366:47]
  wire [6:0] _T_1651 = {io_in_bits_DecodeIn_data_src2[5],_GEN_360}; // @[Cat.scala 30:58]
  wire [5:0] _T_1666 = {io_in_bits_DecodeIn_data_src2[4],io_in_bits_DecodeIn_data_src2[4:0]}; // @[Cat.scala 30:58]
  wire [6:0] _T_1667 = io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isLR_32 ? _T_1651 : {{1'd0}, _T_1666}; // @[PALU.scala 517:22]
  wire [63:0] _WIRE_197 = {{57'd0}, _T_1667};
  wire [5:0] _T_1671 = _T_1636 ? _WIRE_197[5:0] : {{1'd0}, _WIRE_197[4:0]}; // @[PALU.scala 518:27]
  wire [63:0] _T_1675 = {32'h0,io_in_bits_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1676 = io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isLs_Q31 ? _T_1675 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 520:34]
  wire  _T_1681 = io_in_bits_Pctrl_isSRAIWU | io_in_bits_Pctrl_isRs_32 | (io_in_bits_Pctrl_isLR_32 |
    io_in_bits_Pctrl_isLR_Q31) & _WIRE_197[6]; // @[PALU.scala 520:130]
  wire [5:0] _T_1685 = _T_1671 - 6'h1; // @[PALU.scala 327:50]
  wire [5:0] _GEN_365 = io_in_bits_Pctrl_Round ? _T_1685 : _T_1671; // @[PALU.scala 327:{32,42}]
  wire [31:0] _T_1686 = _T_1676[31:0]; // @[PALU.scala 329:42]
  wire [31:0] _T_1688 = $signed(_T_1686) >>> _GEN_365; // @[PALU.scala 329:62]
  wire [31:0] _T_1689 = _T_1676[31:0] >> _GEN_365; // @[PALU.scala 331:41]
  wire [31:0] _GEN_366 = io_in_bits_Pctrl_Arithmetic ? _T_1688 : _T_1689; // @[PALU.scala 328:37 329:29 331:29]
  wire [32:0] _T_1691 = {_GEN_366[31],_GEN_366}; // @[Cat.scala 30:58]
  wire [32:0] _T_1692 = {1'h0,_GEN_366}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_367 = io_in_bits_Pctrl_Arithmetic ? _T_1691 : _T_1692; // @[PALU.scala 96:24 97:15 99:15]
  wire [32:0] _T_1694 = _GEN_367 + 33'h1; // @[PALU.scala 334:66]
  wire [31:0] _GEN_368 = io_in_bits_Pctrl_Round ? _T_1694[32:1] : _GEN_366; // @[PALU.scala 333:32 334:29 336:29]
  wire [31:0] _T_1705 = _T_1676[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1706 = {_T_1705,_T_1676[31:0]}; // @[Cat.scala 30:58]
  wire [126:0] _GEN_49 = {{63'd0}, _T_1706}; // @[PALU.scala 341:35]
  wire [126:0] _T_1707 = _GEN_49 << _T_1671; // @[PALU.scala 341:35]
  wire [126:0] _T_1712 = 127'hffffffffffffffff ^ _T_1707; // @[PALU.scala 345:80]
  wire [126:0] _GEN_369 = _T_1707[63] ? _T_1712 : _T_1707; // @[PALU.scala 345:{53,59}]
  wire  _T_1714 = _GEN_369[63:31] != 33'h0; // @[PALU.scala 346:54]
  wire [31:0] _GEN_370 = _T_1707[63] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 348:57 349:37 351:37]
  wire [31:0] _GEN_372 = _GEN_369[63:31] != 33'h0 ? _GEN_370 : _T_1707[31:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_373 = io_in_bits_Pctrl_ShiftSigned & _T_1714; // @[PALU.scala 343:38 317:45]
  wire [31:0] _GEN_374 = io_in_bits_Pctrl_ShiftSigned ? _GEN_372 : _T_1707[31:0]; // @[PALU.scala 342:25 343:38]
  wire [31:0] _GEN_375 = _T_1681 ? _GEN_368 : _GEN_374; // @[PALU.scala 323:32]
  wire  _GEN_376 = _T_1681 ? 1'h0 : _GEN_373; // @[PALU.scala 323:32 317:45]
  wire [31:0] _GEN_377 = _T_1671 != 6'h0 ? _GEN_375 : _T_1676[31:0]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_378 = _T_1671 != 6'h0 & _GEN_376; // @[PALU.scala 322:31 317:45]
  wire [31:0] _T_1740 = _T_1676[63:32]; // @[PALU.scala 329:42]
  wire [31:0] _T_1742 = $signed(_T_1740) >>> _GEN_365; // @[PALU.scala 329:62]
  wire [31:0] _T_1743 = _T_1676[63:32] >> _GEN_365; // @[PALU.scala 331:41]
  wire [31:0] _GEN_380 = io_in_bits_Pctrl_Arithmetic ? _T_1742 : _T_1743; // @[PALU.scala 328:37 329:29 331:29]
  wire [32:0] _T_1745 = {_GEN_380[31],_GEN_380}; // @[Cat.scala 30:58]
  wire [32:0] _T_1746 = {1'h0,_GEN_380}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_381 = io_in_bits_Pctrl_Arithmetic ? _T_1745 : _T_1746; // @[PALU.scala 96:24 97:15 99:15]
  wire [32:0] _T_1748 = _GEN_381 + 33'h1; // @[PALU.scala 334:66]
  wire [31:0] _GEN_382 = io_in_bits_Pctrl_Round ? _T_1748[32:1] : _GEN_380; // @[PALU.scala 333:32 334:29 336:29]
  wire [31:0] _T_1759 = _T_1676[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1760 = {_T_1759,_T_1676[63:32]}; // @[Cat.scala 30:58]
  wire [126:0] _GEN_52 = {{63'd0}, _T_1760}; // @[PALU.scala 341:35]
  wire [126:0] _T_1761 = _GEN_52 << _T_1671; // @[PALU.scala 341:35]
  wire [126:0] _T_1766 = 127'hffffffffffffffff ^ _T_1761; // @[PALU.scala 345:80]
  wire [126:0] _GEN_383 = _T_1761[63] ? _T_1766 : _T_1761; // @[PALU.scala 345:{53,59}]
  wire  _T_1768 = _GEN_383[63:31] != 33'h0; // @[PALU.scala 346:54]
  wire [31:0] _GEN_384 = _T_1761[63] ? 32'h80000000 : 32'h7fffffff; // @[PALU.scala 348:57 349:37 351:37]
  wire [31:0] _GEN_386 = _GEN_383[63:31] != 33'h0 ? _GEN_384 : _T_1761[31:0]; // @[PALU.scala 342:25 346:62]
  wire  _GEN_387 = io_in_bits_Pctrl_ShiftSigned & _T_1768; // @[PALU.scala 343:38 317:45]
  wire [31:0] _GEN_388 = io_in_bits_Pctrl_ShiftSigned ? _GEN_386 : _T_1761[31:0]; // @[PALU.scala 342:25 343:38]
  wire [31:0] _GEN_389 = _T_1681 ? _GEN_382 : _GEN_388; // @[PALU.scala 323:32]
  wire  _GEN_390 = _T_1681 ? 1'h0 : _GEN_387; // @[PALU.scala 323:32 317:45]
  wire [31:0] _GEN_391 = _T_1671 != 6'h0 ? _GEN_389 : _T_1676[63:32]; // @[PALU.scala 321:17 322:31]
  wire  _GEN_392 = _T_1671 != 6'h0 & _GEN_390; // @[PALU.scala 322:31 317:45]
  wire  _T_1790 = _GEN_378 | _GEN_392; // @[PALU.scala 361:24]
  wire [64:0] _T_1792 = {_T_1790,_GEN_391,_GEN_377}; // @[Cat.scala 30:58]
  wire [31:0] _T_1798 = _T_1792[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1799 = {_T_1798,_T_1792[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1801 = io_in_bits_Pctrl_isLs_Q31 | io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isSRAIWU ? _T_1799 :
    _T_1792[63:0]; // @[PALU.scala 521:26]
  wire [6:0] _T_1827 = {io_in_bits_DecodeIn_data_src2[5],io_in_bits_DecodeIn_data_src2[5:0]}; // @[Cat.scala 30:58]
  wire [5:0] _T_1830 = io_in_bits_Pctrl_isRs_XLEN ? _T_1827[5:0] : {{1'd0}, _T_1827[4:0]}; // @[PALU.scala 526:27]
  wire [63:0] _T_1835 = {io_in_bits_DecodeIn_data_src1[31:0],io_in_bits_DecodeIn_data_src3[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1838 = {io_in_bits_DecodeIn_data_src3[31:0],io_in_bits_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1839 = _T_1827[5] ? _T_1835 : _T_1838; // @[PALU.scala 527:47]
  wire [63:0] _T_1840 = io_in_bits_Pctrl_isFSRW ? _T_1839 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 527:36]
  wire  _T_1841 = io_in_bits_Pctrl_isRs_XLEN & io_in_bits_Pctrl_Round; // @[PALU.scala 527:144]
  wire  _T_1843 = io_in_bits_Pctrl_isRs_XLEN & io_in_bits_Pctrl_Arithmetic; // @[PALU.scala 527:215]
  wire [5:0] _T_1847 = _T_1830 - 6'h1; // @[PALU.scala 327:50]
  wire [5:0] _GEN_396 = _T_1841 ? _T_1847 : _T_1830; // @[PALU.scala 327:{32,42}]
  wire [63:0] _T_1848 = io_in_bits_Pctrl_isFSRW ? _T_1839 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 329:42]
  wire [63:0] _T_1850 = $signed(_T_1848) >>> _GEN_396; // @[PALU.scala 329:62]
  wire [63:0] _T_1851 = _T_1840 >> _GEN_396; // @[PALU.scala 331:41]
  wire [63:0] _GEN_397 = _T_1843 ? _T_1850 : _T_1851; // @[PALU.scala 328:37 329:29 331:29]
  wire [64:0] _T_1853 = {_GEN_397[63],_GEN_397}; // @[Cat.scala 30:58]
  wire [64:0] _T_1854 = {1'h0,_GEN_397}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_398 = _T_1843 ? _T_1853 : _T_1854; // @[PALU.scala 96:24 97:15 99:15]
  wire [64:0] _T_1856 = _GEN_398 + 65'h1; // @[PALU.scala 334:66]
  wire [63:0] _GEN_399 = _T_1841 ? _T_1856[64:1] : _GEN_397; // @[PALU.scala 333:32 334:29 336:29]
  wire [63:0] _GEN_408 = _T_1830 != 6'h0 ? _GEN_399 : _T_1840; // @[PALU.scala 321:17 322:31]
  wire [64:0] _T_1898 = {1'h0,_GEN_408}; // @[Cat.scala 30:58]
  wire [31:0] _T_1903 = _T_1898[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1904 = {_T_1903,_T_1898[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_1905 = io_in_bits_Pctrl_isRs_XLEN ? _T_1898[63:0] : _T_1904; // @[PALU.scala 528:26]
  wire [63:0] _GEN_410 = io_in_bits_Pctrl_isRs_XLEN | io_in_bits_Pctrl_isFSRW | io_in_bits_Pctrl_isWext ? _T_1905 :
    io_in_bits_DecodeIn_data_src1; // @[PALU.scala 524:44 528:20]
  wire  _GEN_411 = (io_in_bits_Pctrl_isRs_XLEN | io_in_bits_Pctrl_isFSRW | io_in_bits_Pctrl_isWext) & _T_1898[64]; // @[PALU.scala 524:44 529:20]
  wire [63:0] _GEN_412 = io_in_bits_Pctrl_isRs_32 | io_in_bits_Pctrl_isLs_32 | io_in_bits_Pctrl_isLR_32 |
    io_in_bits_Pctrl_isLs_Q31 | io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isSRAIWU ? _T_1801 : _GEN_410; // @[PALU.scala 515:77 521:20]
  wire  _GEN_413 = io_in_bits_Pctrl_isRs_32 | io_in_bits_Pctrl_isLs_32 | io_in_bits_Pctrl_isLR_32 |
    io_in_bits_Pctrl_isLs_Q31 | io_in_bits_Pctrl_isLR_Q31 | io_in_bits_Pctrl_isSRAIWU ? _T_1792[64] : _GEN_411; // @[PALU.scala 515:77 522:20]
  wire [63:0] _GEN_414 = io_in_bits_Pctrl_isRs_8 | io_in_bits_Pctrl_isLs_8 | io_in_bits_Pctrl_isLR_8 ? _T_1620[63:0] :
    _GEN_412; // @[PALU.scala 506:40 512:20]
  wire  _GEN_415 = io_in_bits_Pctrl_isRs_8 | io_in_bits_Pctrl_isLs_8 | io_in_bits_Pctrl_isLR_8 ? _T_1620[64] : _GEN_413; // @[PALU.scala 506:40 513:20]
  wire [63:0] shifterRes = io_in_bits_Pctrl_isRs_16 | io_in_bits_Pctrl_isLs_16 | io_in_bits_Pctrl_isLR_16 ? _T_1130[63:0
    ] : _GEN_414; // @[PALU.scala 498:37 504:20]
  wire  shifterOV = io_in_bits_Pctrl_isRs_16 | io_in_bits_Pctrl_isLs_16 | io_in_bits_Pctrl_isLR_16 ? _T_1130[64] :
    _GEN_415; // @[PALU.scala 498:37 505:20]
  wire  _T_1909 = ~io_in_bits_DecodeIn_ctrl_func24; // @[PALU.scala 534:44]
  wire [15:0] _T_1914 = io_in_bits_DecodeIn_data_src1[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1916 = _T_1914 ^ io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_418 = _T_1909 ? _T_1916 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_1918 = _GEN_418 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire [30:0] _T_1920 = 31'hffff << io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 389:46]
  wire  _T_1921 = _T_1918 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_1925 = 16'hffff ^ _T_1920[15:0]; // @[PALU.scala 392:76]
  wire [15:0] _T_1926 = io_in_bits_DecodeIn_data_src1[15] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_1929 = ~_T_1909 & _T_1921; // @[PALU.scala 393:36]
  wire [15:0] _T_1933 = io_in_bits_DecodeIn_data_src1[15] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_420 = ~_T_1909 & _T_1921 ? _T_1933 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_421 = _T_1918 != 16'h0 & _T_1909 | _T_1929; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_422 = _T_1918 != 16'h0 & _T_1909 ? _T_1926 : _GEN_420; // @[PALU.scala 390:44 392:21]
  wire [15:0] _T_1945 = io_in_bits_DecodeIn_data_src1[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1947 = _T_1945 ^ io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_423 = _T_1909 ? _T_1947 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_1949 = _GEN_423 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire  _T_1952 = _T_1949 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_1957 = io_in_bits_DecodeIn_data_src1[31] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_1960 = ~_T_1909 & _T_1952; // @[PALU.scala 393:36]
  wire [15:0] _T_1964 = io_in_bits_DecodeIn_data_src1[31] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_425 = ~_T_1909 & _T_1952 ? _T_1964 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_426 = _T_1949 != 16'h0 & _T_1909 | _T_1960; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_427 = _T_1949 != 16'h0 & _T_1909 ? _T_1957 : _GEN_425; // @[PALU.scala 390:44 392:21]
  wire [15:0] _T_1976 = io_in_bits_DecodeIn_data_src1[47] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_1978 = _T_1976 ^ io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_428 = _T_1909 ? _T_1978 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_1980 = _GEN_428 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire  _T_1983 = _T_1980 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_1988 = io_in_bits_DecodeIn_data_src1[47] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_1991 = ~_T_1909 & _T_1983; // @[PALU.scala 393:36]
  wire [15:0] _T_1995 = io_in_bits_DecodeIn_data_src1[47] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_430 = ~_T_1909 & _T_1983 ? _T_1995 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_431 = _T_1980 != 16'h0 & _T_1909 | _T_1991; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_432 = _T_1980 != 16'h0 & _T_1909 ? _T_1988 : _GEN_430; // @[PALU.scala 390:44 392:21]
  wire [15:0] _T_2007 = io_in_bits_DecodeIn_data_src1[63] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2009 = _T_2007 ^ io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 384:58]
  wire [15:0] _GEN_433 = _T_1909 ? _T_2009 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 383:29 384:22 386:22]
  wire [15:0] _T_2011 = _GEN_433 >> io_in_bits_DecodeIn_data_src2[3:0]; // @[PALU.scala 388:28]
  wire  _T_2014 = _T_2011 != 16'h0; // @[PALU.scala 390:22]
  wire [15:0] _T_2019 = io_in_bits_DecodeIn_data_src1[63] ? _T_1920[15:0] : _T_1925; // @[PALU.scala 392:27]
  wire  _T_2022 = ~_T_1909 & _T_2014; // @[PALU.scala 393:36]
  wire [15:0] _T_2026 = io_in_bits_DecodeIn_data_src1[63] ? 16'h0 : _T_1925; // @[PALU.scala 395:27]
  wire [15:0] _GEN_435 = ~_T_1909 & _T_2014 ? _T_2026 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_436 = _T_2011 != 16'h0 & _T_1909 | _T_2022; // @[PALU.scala 390:44 391:23]
  wire [15:0] _GEN_437 = _T_2011 != 16'h0 & _T_1909 ? _T_2019 : _GEN_435; // @[PALU.scala 390:44 392:21]
  wire  _T_2036 = _GEN_421 | _GEN_426 | _GEN_431 | _GEN_436; // @[PALU.scala 400:24]
  wire [64:0] _T_2040 = {_T_2036,_GEN_437,_GEN_432,_GEN_427,_GEN_422}; // @[Cat.scala 30:58]
  wire [7:0] _T_2049 = io_in_bits_DecodeIn_data_src1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2051 = _T_2049 ^ io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_438 = _T_1909 ? _T_2051 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2053 = _GEN_438 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire [14:0] _T_2055 = 15'hff << io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 389:46]
  wire  _T_2056 = _T_2053 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2060 = 8'hff ^ _T_2055[7:0]; // @[PALU.scala 392:76]
  wire [7:0] _T_2061 = io_in_bits_DecodeIn_data_src1[7] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2064 = ~_T_1909 & _T_2056; // @[PALU.scala 393:36]
  wire [7:0] _T_2068 = io_in_bits_DecodeIn_data_src1[7] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_440 = ~_T_1909 & _T_2056 ? _T_2068 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_441 = _T_2053 != 8'h0 & _T_1909 | _T_2064; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_442 = _T_2053 != 8'h0 & _T_1909 ? _T_2061 : _GEN_440; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2080 = io_in_bits_DecodeIn_data_src1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2082 = _T_2080 ^ io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_443 = _T_1909 ? _T_2082 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2084 = _GEN_443 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2087 = _T_2084 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2092 = io_in_bits_DecodeIn_data_src1[15] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2095 = ~_T_1909 & _T_2087; // @[PALU.scala 393:36]
  wire [7:0] _T_2099 = io_in_bits_DecodeIn_data_src1[15] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_445 = ~_T_1909 & _T_2087 ? _T_2099 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_446 = _T_2084 != 8'h0 & _T_1909 | _T_2095; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_447 = _T_2084 != 8'h0 & _T_1909 ? _T_2092 : _GEN_445; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2111 = io_in_bits_DecodeIn_data_src1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2113 = _T_2111 ^ io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_448 = _T_1909 ? _T_2113 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2115 = _GEN_448 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2118 = _T_2115 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2123 = io_in_bits_DecodeIn_data_src1[23] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2126 = ~_T_1909 & _T_2118; // @[PALU.scala 393:36]
  wire [7:0] _T_2130 = io_in_bits_DecodeIn_data_src1[23] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_450 = ~_T_1909 & _T_2118 ? _T_2130 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_451 = _T_2115 != 8'h0 & _T_1909 | _T_2126; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_452 = _T_2115 != 8'h0 & _T_1909 ? _T_2123 : _GEN_450; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2142 = io_in_bits_DecodeIn_data_src1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2144 = _T_2142 ^ io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_453 = _T_1909 ? _T_2144 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2146 = _GEN_453 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2149 = _T_2146 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2154 = io_in_bits_DecodeIn_data_src1[31] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2157 = ~_T_1909 & _T_2149; // @[PALU.scala 393:36]
  wire [7:0] _T_2161 = io_in_bits_DecodeIn_data_src1[31] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_455 = ~_T_1909 & _T_2149 ? _T_2161 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_456 = _T_2146 != 8'h0 & _T_1909 | _T_2157; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_457 = _T_2146 != 8'h0 & _T_1909 ? _T_2154 : _GEN_455; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2173 = io_in_bits_DecodeIn_data_src1[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2175 = _T_2173 ^ io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_458 = _T_1909 ? _T_2175 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2177 = _GEN_458 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2180 = _T_2177 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2185 = io_in_bits_DecodeIn_data_src1[39] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2188 = ~_T_1909 & _T_2180; // @[PALU.scala 393:36]
  wire [7:0] _T_2192 = io_in_bits_DecodeIn_data_src1[39] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_460 = ~_T_1909 & _T_2180 ? _T_2192 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_461 = _T_2177 != 8'h0 & _T_1909 | _T_2188; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_462 = _T_2177 != 8'h0 & _T_1909 ? _T_2185 : _GEN_460; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2204 = io_in_bits_DecodeIn_data_src1[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2206 = _T_2204 ^ io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_463 = _T_1909 ? _T_2206 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2208 = _GEN_463 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2211 = _T_2208 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2216 = io_in_bits_DecodeIn_data_src1[47] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2219 = ~_T_1909 & _T_2211; // @[PALU.scala 393:36]
  wire [7:0] _T_2223 = io_in_bits_DecodeIn_data_src1[47] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_465 = ~_T_1909 & _T_2211 ? _T_2223 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_466 = _T_2208 != 8'h0 & _T_1909 | _T_2219; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_467 = _T_2208 != 8'h0 & _T_1909 ? _T_2216 : _GEN_465; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2235 = io_in_bits_DecodeIn_data_src1[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2237 = _T_2235 ^ io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_468 = _T_1909 ? _T_2237 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2239 = _GEN_468 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2242 = _T_2239 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2247 = io_in_bits_DecodeIn_data_src1[55] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2250 = ~_T_1909 & _T_2242; // @[PALU.scala 393:36]
  wire [7:0] _T_2254 = io_in_bits_DecodeIn_data_src1[55] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_470 = ~_T_1909 & _T_2242 ? _T_2254 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_471 = _T_2239 != 8'h0 & _T_1909 | _T_2250; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_472 = _T_2239 != 8'h0 & _T_1909 ? _T_2247 : _GEN_470; // @[PALU.scala 390:44 392:21]
  wire [7:0] _T_2266 = io_in_bits_DecodeIn_data_src1[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2268 = _T_2266 ^ io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 384:58]
  wire [7:0] _GEN_473 = _T_1909 ? _T_2268 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 383:29 384:22 386:22]
  wire [7:0] _T_2270 = _GEN_473 >> io_in_bits_DecodeIn_data_src2[2:0]; // @[PALU.scala 388:28]
  wire  _T_2273 = _T_2270 != 8'h0; // @[PALU.scala 390:22]
  wire [7:0] _T_2278 = io_in_bits_DecodeIn_data_src1[63] ? _T_2055[7:0] : _T_2060; // @[PALU.scala 392:27]
  wire  _T_2281 = ~_T_1909 & _T_2273; // @[PALU.scala 393:36]
  wire [7:0] _T_2285 = io_in_bits_DecodeIn_data_src1[63] ? 8'h0 : _T_2060; // @[PALU.scala 395:27]
  wire [7:0] _GEN_475 = ~_T_1909 & _T_2273 ? _T_2285 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_476 = _T_2270 != 8'h0 & _T_1909 | _T_2281; // @[PALU.scala 390:44 391:23]
  wire [7:0] _GEN_477 = _T_2270 != 8'h0 & _T_1909 ? _T_2278 : _GEN_475; // @[PALU.scala 390:44 392:21]
  wire  _T_2299 = _GEN_441 | _GEN_446 | _GEN_451 | _GEN_456 | _GEN_461 | _GEN_466 | _GEN_471 | _GEN_476; // @[PALU.scala 400:24]
  wire [64:0] _T_2307 = {_T_2299,_GEN_477,_GEN_472,_GEN_467,_GEN_462,_GEN_457,_GEN_452,_GEN_447,_GEN_442}; // @[Cat.scala 30:58]
  wire [31:0] _T_2317 = io_in_bits_DecodeIn_data_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2319 = _T_2317 ^ io_in_bits_DecodeIn_data_src1[31:0]; // @[PALU.scala 384:58]
  wire [31:0] _GEN_478 = _T_15 ? _T_2319 : io_in_bits_DecodeIn_data_src1[31:0]; // @[PALU.scala 383:29 384:22 386:22]
  wire [31:0] _T_2321 = _GEN_478 >> io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 388:28]
  wire [62:0] _T_2323 = 63'hffffffff << io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 389:46]
  wire  _T_2324 = _T_2321 != 32'h0; // @[PALU.scala 390:22]
  wire [31:0] _T_2328 = 32'hffffffff ^ _T_2323[31:0]; // @[PALU.scala 392:76]
  wire [31:0] _T_2329 = io_in_bits_DecodeIn_data_src1[31] ? _T_2323[31:0] : _T_2328; // @[PALU.scala 392:27]
  wire  _T_2332 = ~_T_15 & _T_2324; // @[PALU.scala 393:36]
  wire [31:0] _T_2336 = io_in_bits_DecodeIn_data_src1[31] ? 32'h0 : _T_2328; // @[PALU.scala 395:27]
  wire [31:0] _GEN_480 = ~_T_15 & _T_2324 ? _T_2336 : io_in_bits_DecodeIn_data_src1[31:0]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_481 = _T_2321 != 32'h0 & _T_15 | _T_2332; // @[PALU.scala 390:44 391:23]
  wire [31:0] _GEN_482 = _T_2321 != 32'h0 & _T_15 ? _T_2329 : _GEN_480; // @[PALU.scala 390:44 392:21]
  wire [31:0] _T_2348 = io_in_bits_DecodeIn_data_src1[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2350 = _T_2348 ^ io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 384:58]
  wire [31:0] _GEN_483 = _T_15 ? _T_2350 : io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 383:29 384:22 386:22]
  wire [31:0] _T_2352 = _GEN_483 >> io_in_bits_DecodeIn_data_src2[4:0]; // @[PALU.scala 388:28]
  wire  _T_2355 = _T_2352 != 32'h0; // @[PALU.scala 390:22]
  wire [31:0] _T_2360 = io_in_bits_DecodeIn_data_src1[63] ? _T_2323[31:0] : _T_2328; // @[PALU.scala 392:27]
  wire  _T_2363 = ~_T_15 & _T_2355; // @[PALU.scala 393:36]
  wire [31:0] _T_2367 = io_in_bits_DecodeIn_data_src1[63] ? 32'h0 : _T_2328; // @[PALU.scala 395:27]
  wire [31:0] _GEN_485 = ~_T_15 & _T_2355 ? _T_2367 : io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 393:51 395:21]
  wire  _GEN_486 = _T_2352 != 32'h0 & _T_15 | _T_2363; // @[PALU.scala 390:44 391:23]
  wire [31:0] _GEN_487 = _T_2352 != 32'h0 & _T_15 ? _T_2360 : _GEN_485; // @[PALU.scala 390:44 392:21]
  wire  _T_2375 = _GEN_481 | _GEN_486; // @[PALU.scala 400:24]
  wire [64:0] _T_2377 = {_T_2375,_GEN_487,_GEN_482}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_488 = io_in_bits_Pctrl_isclip_32 ? _T_2377[63:0] : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 541:26 543:17]
  wire  _GEN_489 = io_in_bits_Pctrl_isclip_32 & _T_2377[64]; // @[PALU.scala 541:26 544:17]
  wire [63:0] _GEN_490 = io_in_bits_Pctrl_isClip_8 ? _T_2307[63:0] : _GEN_488; // @[PALU.scala 537:25 539:17]
  wire  _GEN_491 = io_in_bits_Pctrl_isClip_8 ? _T_2307[64] : _GEN_489; // @[PALU.scala 537:25 540:17]
  wire [63:0] clipRes = io_in_bits_Pctrl_isClip_16 ? _T_2040[63:0] : _GEN_490; // @[PALU.scala 533:20 535:17]
  wire  clipOV = io_in_bits_Pctrl_isClip_16 ? _T_2040[64] : _GEN_491; // @[PALU.scala 533:20 536:17]
  wire  _T_2384 = io_in_bits_DecodeIn_data_src1[15:0] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2390 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 413:42]
  wire [15:0] _T_2392 = _T_2390 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_494 = io_in_bits_DecodeIn_data_src1[15] ? _T_2392 : io_in_bits_DecodeIn_data_src1[15:0]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_496 = io_in_bits_DecodeIn_data_src1[15:0] == 16'h8000 ? 16'h7fff : _GEN_494; // @[PALU.scala 409:53 411:23]
  wire  _T_2397 = io_in_bits_DecodeIn_data_src1[31:16] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2403 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 413:42]
  wire [15:0] _T_2405 = _T_2403 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_497 = io_in_bits_DecodeIn_data_src1[31] ? _T_2405 : io_in_bits_DecodeIn_data_src1[31:16]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_499 = io_in_bits_DecodeIn_data_src1[31:16] == 16'h8000 ? 16'h7fff : _GEN_497; // @[PALU.scala 409:53 411:23]
  wire  _T_2410 = io_in_bits_DecodeIn_data_src1[47:32] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2416 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 413:42]
  wire [15:0] _T_2418 = _T_2416 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_500 = io_in_bits_DecodeIn_data_src1[47] ? _T_2418 : io_in_bits_DecodeIn_data_src1[47:32]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_502 = io_in_bits_DecodeIn_data_src1[47:32] == 16'h8000 ? 16'h7fff : _GEN_500; // @[PALU.scala 409:53 411:23]
  wire  _T_2423 = io_in_bits_DecodeIn_data_src1[63:48] == 16'h8000; // @[PALU.scala 409:22]
  wire [15:0] _T_2429 = 16'hffff ^ io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 413:42]
  wire [15:0] _T_2431 = _T_2429 + 16'h1; // @[PALU.scala 413:48]
  wire [15:0] _GEN_503 = io_in_bits_DecodeIn_data_src1[63] ? _T_2431 : io_in_bits_DecodeIn_data_src1[63:48]; // @[PALU.scala 412:44 413:23]
  wire [15:0] _GEN_505 = io_in_bits_DecodeIn_data_src1[63:48] == 16'h8000 ? 16'h7fff : _GEN_503; // @[PALU.scala 409:53 411:23]
  wire  _T_2434 = _T_2384 | _T_2397 | _T_2410 | _T_2423; // @[PALU.scala 417:24]
  wire [64:0] _T_2438 = {_T_2434,_GEN_505,_GEN_502,_GEN_499,_GEN_496}; // @[Cat.scala 30:58]
  wire  _T_2445 = io_in_bits_DecodeIn_data_src1[7:0] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2451 = 8'hff ^ io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 413:42]
  wire [7:0] _T_2453 = _T_2451 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_506 = io_in_bits_DecodeIn_data_src1[7] ? _T_2453 : io_in_bits_DecodeIn_data_src1[7:0]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_508 = io_in_bits_DecodeIn_data_src1[7:0] == 8'h80 ? 8'h7f : _GEN_506; // @[PALU.scala 409:53 411:23]
  wire  _T_2458 = io_in_bits_DecodeIn_data_src1[15:8] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2464 = 8'hff ^ io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 413:42]
  wire [7:0] _T_2466 = _T_2464 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_509 = io_in_bits_DecodeIn_data_src1[15] ? _T_2466 : io_in_bits_DecodeIn_data_src1[15:8]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_511 = io_in_bits_DecodeIn_data_src1[15:8] == 8'h80 ? 8'h7f : _GEN_509; // @[PALU.scala 409:53 411:23]
  wire  _T_2471 = io_in_bits_DecodeIn_data_src1[23:16] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2477 = 8'hff ^ io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 413:42]
  wire [7:0] _T_2479 = _T_2477 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_512 = io_in_bits_DecodeIn_data_src1[23] ? _T_2479 : io_in_bits_DecodeIn_data_src1[23:16]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_514 = io_in_bits_DecodeIn_data_src1[23:16] == 8'h80 ? 8'h7f : _GEN_512; // @[PALU.scala 409:53 411:23]
  wire  _T_2484 = io_in_bits_DecodeIn_data_src1[31:24] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2490 = 8'hff ^ io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 413:42]
  wire [7:0] _T_2492 = _T_2490 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_515 = io_in_bits_DecodeIn_data_src1[31] ? _T_2492 : io_in_bits_DecodeIn_data_src1[31:24]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_517 = io_in_bits_DecodeIn_data_src1[31:24] == 8'h80 ? 8'h7f : _GEN_515; // @[PALU.scala 409:53 411:23]
  wire  _T_2497 = io_in_bits_DecodeIn_data_src1[39:32] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2503 = 8'hff ^ io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 413:42]
  wire [7:0] _T_2505 = _T_2503 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_518 = io_in_bits_DecodeIn_data_src1[39] ? _T_2505 : io_in_bits_DecodeIn_data_src1[39:32]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_520 = io_in_bits_DecodeIn_data_src1[39:32] == 8'h80 ? 8'h7f : _GEN_518; // @[PALU.scala 409:53 411:23]
  wire  _T_2510 = io_in_bits_DecodeIn_data_src1[47:40] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2516 = 8'hff ^ io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 413:42]
  wire [7:0] _T_2518 = _T_2516 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_521 = io_in_bits_DecodeIn_data_src1[47] ? _T_2518 : io_in_bits_DecodeIn_data_src1[47:40]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_523 = io_in_bits_DecodeIn_data_src1[47:40] == 8'h80 ? 8'h7f : _GEN_521; // @[PALU.scala 409:53 411:23]
  wire  _T_2523 = io_in_bits_DecodeIn_data_src1[55:48] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2529 = 8'hff ^ io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 413:42]
  wire [7:0] _T_2531 = _T_2529 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_524 = io_in_bits_DecodeIn_data_src1[55] ? _T_2531 : io_in_bits_DecodeIn_data_src1[55:48]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_526 = io_in_bits_DecodeIn_data_src1[55:48] == 8'h80 ? 8'h7f : _GEN_524; // @[PALU.scala 409:53 411:23]
  wire  _T_2536 = io_in_bits_DecodeIn_data_src1[63:56] == 8'h80; // @[PALU.scala 409:22]
  wire [7:0] _T_2542 = 8'hff ^ io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 413:42]
  wire [7:0] _T_2544 = _T_2542 + 8'h1; // @[PALU.scala 413:48]
  wire [7:0] _GEN_527 = io_in_bits_DecodeIn_data_src1[63] ? _T_2544 : io_in_bits_DecodeIn_data_src1[63:56]; // @[PALU.scala 412:44 413:23]
  wire [7:0] _GEN_529 = io_in_bits_DecodeIn_data_src1[63:56] == 8'h80 ? 8'h7f : _GEN_527; // @[PALU.scala 409:53 411:23]
  wire  _T_2551 = _T_2445 | _T_2458 | _T_2471 | _T_2484 | _T_2497 | _T_2510 | _T_2523 | _T_2536; // @[PALU.scala 417:24]
  wire [64:0] _T_2559 = {_T_2551,_GEN_529,_GEN_526,_GEN_523,_GEN_520,_GEN_517,_GEN_514,_GEN_511,_GEN_508}; // @[Cat.scala 30:58]
  wire [63:0] _T_2565 = io_in_bits_Pctrl_isSat_W ? _T_1675 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 558:35]
  wire  _T_2570 = _T_2565[31:0] == 32'h80000000; // @[PALU.scala 409:22]
  wire [31:0] _T_2576 = 32'hffffffff ^ _T_2565[31:0]; // @[PALU.scala 413:42]
  wire [31:0] _T_2578 = _T_2576 + 32'h1; // @[PALU.scala 413:48]
  wire [31:0] _GEN_530 = _T_2565[31] ? _T_2578 : _T_2565[31:0]; // @[PALU.scala 412:44 413:23]
  wire [31:0] _GEN_532 = _T_2565[31:0] == 32'h80000000 ? 32'h7fffffff : _GEN_530; // @[PALU.scala 409:53 411:23]
  wire  _T_2583 = _T_2565[63:32] == 32'h80000000; // @[PALU.scala 409:22]
  wire [31:0] _T_2589 = 32'hffffffff ^ _T_2565[63:32]; // @[PALU.scala 413:42]
  wire [31:0] _T_2591 = _T_2589 + 32'h1; // @[PALU.scala 413:48]
  wire [31:0] _GEN_533 = _T_2565[63] ? _T_2591 : _T_2565[63:32]; // @[PALU.scala 412:44 413:23]
  wire [31:0] _GEN_535 = _T_2565[63:32] == 32'h80000000 ? 32'h7fffffff : _GEN_533; // @[PALU.scala 409:53 411:23]
  wire  _T_2592 = _T_2570 | _T_2583; // @[PALU.scala 417:24]
  wire [64:0] _T_2594 = {_T_2592,_GEN_535,_GEN_532}; // @[Cat.scala 30:58]
  wire [31:0] _T_2598 = _T_2594[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2599 = {_T_2598,_T_2594[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2601 = io_in_bits_Pctrl_isSat_W ? _T_2599 : _T_2594[63:0]; // @[PALU.scala 559:22]
  wire [63:0] _GEN_536 = io_in_bits_Pctrl_isSat_32 | io_in_bits_Pctrl_isSat_W ? _T_2601 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 557:35 559:16]
  wire  _GEN_537 = (io_in_bits_Pctrl_isSat_32 | io_in_bits_Pctrl_isSat_W) & _T_2594[64]; // @[PALU.scala 557:35 560:16]
  wire [63:0] _GEN_538 = io_in_bits_Pctrl_isSat_8 ? _T_2559[63:0] : _GEN_536; // @[PALU.scala 553:24 555:16]
  wire  _GEN_539 = io_in_bits_Pctrl_isSat_8 ? _T_2559[64] : _GEN_537; // @[PALU.scala 553:24 556:16]
  wire [63:0] satRes = io_in_bits_Pctrl_isSat_16 ? _T_2438[63:0] : _GEN_538; // @[PALU.scala 549:19 551:16]
  wire  satOV = io_in_bits_Pctrl_isSat_16 ? _T_2438[64] : _GEN_539; // @[PALU.scala 549:19 552:16]
  wire [4:0] _T_2604 = io_in_bits_DecodeIn_data_src2[4:0] & 5'h1b; // @[PALU.scala 566:45]
  wire  _T_2607 = ~io_in_bits_DecodeIn_data_src2[2]; // @[PALU.scala 566:57]
  wire [7:0] _T_2616 = io_in_bits_DecodeIn_data_src1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2617 = {_T_2616,io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2618 = {8'h0,io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_542 = _T_2607 ? _T_2617 : _T_2618; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2626 = io_in_bits_DecodeIn_data_src1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2627 = {_T_2626,io_in_bits_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2628 = {8'h0,io_in_bits_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_543 = _T_2607 ? _T_2627 : _T_2628; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2635 = io_in_bits_DecodeIn_data_src1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2636 = {_T_2635,io_in_bits_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2637 = {8'h0,io_in_bits_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_544 = _T_2607 ? _T_2636 : _T_2637; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2638 = _T_2604 == 5'h9 ? _GEN_543 : _GEN_544; // @[PALU.scala 464:107]
  wire [15:0] _T_2639 = _T_2604 == 5'h8 ? _GEN_542 : _T_2638; // @[PALU.scala 464:26]
  wire [7:0] _T_2666 = io_in_bits_DecodeIn_data_src1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2667 = {_T_2666,io_in_bits_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2668 = {8'h0,io_in_bits_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_547 = _T_2607 ? _T_2667 : _T_2668; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2669 = _T_2604 == 5'hb ? _GEN_542 : _GEN_547; // @[PALU.scala 465:107]
  wire [15:0] _T_2670 = _T_2604 == 5'h13 ? _GEN_543 : _T_2669; // @[PALU.scala 465:26]
  wire [7:0] _T_2680 = io_in_bits_DecodeIn_data_src1[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2681 = {_T_2680,io_in_bits_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2682 = {8'h0,io_in_bits_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_548 = _T_2607 ? _T_2681 : _T_2682; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2690 = io_in_bits_DecodeIn_data_src1[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2691 = {_T_2690,io_in_bits_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2692 = {8'h0,io_in_bits_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_549 = _T_2607 ? _T_2691 : _T_2692; // @[PALU.scala 96:24 97:15 99:15]
  wire [7:0] _T_2699 = io_in_bits_DecodeIn_data_src1[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2700 = {_T_2699,io_in_bits_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2701 = {8'h0,io_in_bits_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_550 = _T_2607 ? _T_2700 : _T_2701; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2702 = _T_2604 == 5'h9 ? _GEN_549 : _GEN_550; // @[PALU.scala 464:107]
  wire [15:0] _T_2703 = _T_2604 == 5'h8 ? _GEN_548 : _T_2702; // @[PALU.scala 464:26]
  wire [7:0] _T_2730 = io_in_bits_DecodeIn_data_src1[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2731 = {_T_2730,io_in_bits_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [15:0] _T_2732 = {8'h0,io_in_bits_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_553 = _T_2607 ? _T_2731 : _T_2732; // @[PALU.scala 96:24 97:15 99:15]
  wire [15:0] _T_2733 = _T_2604 == 5'hb ? _GEN_548 : _GEN_553; // @[PALU.scala 465:107]
  wire [15:0] _T_2734 = _T_2604 == 5'h13 ? _GEN_549 : _T_2733; // @[PALU.scala 465:26]
  wire [63:0] _T_2736 = {_T_2703,_T_2734,_T_2639,_T_2670}; // @[Cat.scala 30:58]
  wire [63:0] unpackRes = io_in_bits_Pctrl_isUnpack ? _T_2736 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 565:19 566:19]
  wire  _T_2740 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[15]; // @[PALU.scala 423:29]
  wire  _T_2742 = io_in_bits_DecodeIn_data_src1[0] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2744 = io_in_bits_DecodeIn_data_src1[1] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2746 = io_in_bits_DecodeIn_data_src1[2] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2748 = io_in_bits_DecodeIn_data_src1[3] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2750 = io_in_bits_DecodeIn_data_src1[4] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2752 = io_in_bits_DecodeIn_data_src1[5] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2754 = io_in_bits_DecodeIn_data_src1[6] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2756 = io_in_bits_DecodeIn_data_src1[7] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2758 = io_in_bits_DecodeIn_data_src1[8] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2760 = io_in_bits_DecodeIn_data_src1[9] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2762 = io_in_bits_DecodeIn_data_src1[10] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2764 = io_in_bits_DecodeIn_data_src1[11] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2766 = io_in_bits_DecodeIn_data_src1[12] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2768 = io_in_bits_DecodeIn_data_src1[13] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2770 = io_in_bits_DecodeIn_data_src1[14] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2772 = io_in_bits_DecodeIn_data_src1[15] == _T_2740; // @[PALU.scala 425:59]
  wire  _T_2774 = _T_2770 & _T_2772; // @[PALU.scala 427:113]
  wire  _T_2776 = _T_2768 & (_T_2770 & _T_2772); // @[PALU.scala 427:113]
  wire  _T_2778 = _T_2766 & (_T_2768 & (_T_2770 & _T_2772)); // @[PALU.scala 427:113]
  wire  _T_2780 = _T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))); // @[PALU.scala 427:113]
  wire  _T_2782 = _T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))); // @[PALU.scala 427:113]
  wire  _T_2784 = _T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))))); // @[PALU.scala 427:113]
  wire  _T_2786 = _T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))))); // @[PALU.scala 427:113]
  wire  _T_2788 = _T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))))))); // @[PALU.scala 427:113]
  wire  _T_2790 = _T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 &
    _T_2772)))))))); // @[PALU.scala 427:113]
  wire  _T_2792 = _T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (
    _T_2770 & _T_2772))))))))); // @[PALU.scala 427:113]
  wire  _T_2794 = _T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (
    _T_2768 & (_T_2770 & _T_2772)))))))))); // @[PALU.scala 427:113]
  wire  _T_2796 = _T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (_T_2764 & (
    _T_2766 & (_T_2768 & (_T_2770 & _T_2772))))))))))); // @[PALU.scala 427:113]
  wire  _T_2798 = _T_2746 & (_T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (_T_2762 & (
    _T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))))))))))); // @[PALU.scala 427:113]
  wire  _T_2800 = _T_2744 & (_T_2746 & (_T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (_T_2760 & (
    _T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772))))))))))))); // @[PALU.scala 427:113]
  wire  _T_2802 = _T_2742 & (_T_2744 & (_T_2746 & (_T_2748 & (_T_2750 & (_T_2752 & (_T_2754 & (_T_2756 & (_T_2758 & (
    _T_2760 & (_T_2762 & (_T_2764 & (_T_2766 & (_T_2768 & (_T_2770 & _T_2772)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_2803 = _T_2772 + _T_2774; // @[PALU.scala 428:38]
  wire [1:0] _GEN_655 = {{1'd0}, _T_2776}; // @[PALU.scala 428:38]
  wire [2:0] _T_2804 = _T_2803 + _GEN_655; // @[PALU.scala 428:38]
  wire [2:0] _GEN_656 = {{2'd0}, _T_2778}; // @[PALU.scala 428:38]
  wire [3:0] _T_2805 = _T_2804 + _GEN_656; // @[PALU.scala 428:38]
  wire [3:0] _GEN_657 = {{3'd0}, _T_2780}; // @[PALU.scala 428:38]
  wire [4:0] _T_2806 = _T_2805 + _GEN_657; // @[PALU.scala 428:38]
  wire [4:0] _GEN_658 = {{4'd0}, _T_2782}; // @[PALU.scala 428:38]
  wire [5:0] _T_2807 = _T_2806 + _GEN_658; // @[PALU.scala 428:38]
  wire [5:0] _GEN_659 = {{5'd0}, _T_2784}; // @[PALU.scala 428:38]
  wire [6:0] _T_2808 = _T_2807 + _GEN_659; // @[PALU.scala 428:38]
  wire [6:0] _GEN_660 = {{6'd0}, _T_2786}; // @[PALU.scala 428:38]
  wire [7:0] _T_2809 = _T_2808 + _GEN_660; // @[PALU.scala 428:38]
  wire [7:0] _GEN_661 = {{7'd0}, _T_2788}; // @[PALU.scala 428:38]
  wire [8:0] _T_2810 = _T_2809 + _GEN_661; // @[PALU.scala 428:38]
  wire [8:0] _GEN_662 = {{8'd0}, _T_2790}; // @[PALU.scala 428:38]
  wire [9:0] _T_2811 = _T_2810 + _GEN_662; // @[PALU.scala 428:38]
  wire [9:0] _GEN_663 = {{9'd0}, _T_2792}; // @[PALU.scala 428:38]
  wire [10:0] _T_2812 = _T_2811 + _GEN_663; // @[PALU.scala 428:38]
  wire [10:0] _GEN_664 = {{10'd0}, _T_2794}; // @[PALU.scala 428:38]
  wire [11:0] _T_2813 = _T_2812 + _GEN_664; // @[PALU.scala 428:38]
  wire [11:0] _GEN_665 = {{11'd0}, _T_2796}; // @[PALU.scala 428:38]
  wire [12:0] _T_2814 = _T_2813 + _GEN_665; // @[PALU.scala 428:38]
  wire [12:0] _GEN_666 = {{12'd0}, _T_2798}; // @[PALU.scala 428:38]
  wire [13:0] _T_2815 = _T_2814 + _GEN_666; // @[PALU.scala 428:38]
  wire [13:0] _GEN_667 = {{13'd0}, _T_2800}; // @[PALU.scala 428:38]
  wire [14:0] _T_2816 = _T_2815 + _GEN_667; // @[PALU.scala 428:38]
  wire [14:0] _GEN_668 = {{14'd0}, _T_2802}; // @[PALU.scala 428:38]
  wire [15:0] _T_2817 = _T_2816 + _GEN_668; // @[PALU.scala 428:38]
  wire [15:0] _T_2819 = _T_2817 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_2820 = io_in_bits_DecodeIn_data_src2[0] ? _T_2817 : _T_2819; // @[PALU.scala 429:26]
  wire  _T_2823 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[31]; // @[PALU.scala 423:29]
  wire  _T_2825 = io_in_bits_DecodeIn_data_src1[16] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2827 = io_in_bits_DecodeIn_data_src1[17] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2829 = io_in_bits_DecodeIn_data_src1[18] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2831 = io_in_bits_DecodeIn_data_src1[19] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2833 = io_in_bits_DecodeIn_data_src1[20] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2835 = io_in_bits_DecodeIn_data_src1[21] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2837 = io_in_bits_DecodeIn_data_src1[22] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2839 = io_in_bits_DecodeIn_data_src1[23] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2841 = io_in_bits_DecodeIn_data_src1[24] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2843 = io_in_bits_DecodeIn_data_src1[25] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2845 = io_in_bits_DecodeIn_data_src1[26] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2847 = io_in_bits_DecodeIn_data_src1[27] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2849 = io_in_bits_DecodeIn_data_src1[28] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2851 = io_in_bits_DecodeIn_data_src1[29] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2853 = io_in_bits_DecodeIn_data_src1[30] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2855 = io_in_bits_DecodeIn_data_src1[31] == _T_2823; // @[PALU.scala 425:59]
  wire  _T_2857 = _T_2853 & _T_2855; // @[PALU.scala 427:113]
  wire  _T_2859 = _T_2851 & (_T_2853 & _T_2855); // @[PALU.scala 427:113]
  wire  _T_2861 = _T_2849 & (_T_2851 & (_T_2853 & _T_2855)); // @[PALU.scala 427:113]
  wire  _T_2863 = _T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))); // @[PALU.scala 427:113]
  wire  _T_2865 = _T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))); // @[PALU.scala 427:113]
  wire  _T_2867 = _T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))))); // @[PALU.scala 427:113]
  wire  _T_2869 = _T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))))); // @[PALU.scala 427:113]
  wire  _T_2871 = _T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))))))); // @[PALU.scala 427:113]
  wire  _T_2873 = _T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 &
    _T_2855)))))))); // @[PALU.scala 427:113]
  wire  _T_2875 = _T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (
    _T_2853 & _T_2855))))))))); // @[PALU.scala 427:113]
  wire  _T_2877 = _T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (
    _T_2851 & (_T_2853 & _T_2855)))))))))); // @[PALU.scala 427:113]
  wire  _T_2879 = _T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (_T_2847 & (
    _T_2849 & (_T_2851 & (_T_2853 & _T_2855))))))))))); // @[PALU.scala 427:113]
  wire  _T_2881 = _T_2829 & (_T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (_T_2845 & (
    _T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))))))))))); // @[PALU.scala 427:113]
  wire  _T_2883 = _T_2827 & (_T_2829 & (_T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (_T_2843 & (
    _T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855))))))))))))); // @[PALU.scala 427:113]
  wire  _T_2885 = _T_2825 & (_T_2827 & (_T_2829 & (_T_2831 & (_T_2833 & (_T_2835 & (_T_2837 & (_T_2839 & (_T_2841 & (
    _T_2843 & (_T_2845 & (_T_2847 & (_T_2849 & (_T_2851 & (_T_2853 & _T_2855)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_2886 = _T_2855 + _T_2857; // @[PALU.scala 428:38]
  wire [1:0] _GEN_669 = {{1'd0}, _T_2859}; // @[PALU.scala 428:38]
  wire [2:0] _T_2887 = _T_2886 + _GEN_669; // @[PALU.scala 428:38]
  wire [2:0] _GEN_670 = {{2'd0}, _T_2861}; // @[PALU.scala 428:38]
  wire [3:0] _T_2888 = _T_2887 + _GEN_670; // @[PALU.scala 428:38]
  wire [3:0] _GEN_671 = {{3'd0}, _T_2863}; // @[PALU.scala 428:38]
  wire [4:0] _T_2889 = _T_2888 + _GEN_671; // @[PALU.scala 428:38]
  wire [4:0] _GEN_672 = {{4'd0}, _T_2865}; // @[PALU.scala 428:38]
  wire [5:0] _T_2890 = _T_2889 + _GEN_672; // @[PALU.scala 428:38]
  wire [5:0] _GEN_673 = {{5'd0}, _T_2867}; // @[PALU.scala 428:38]
  wire [6:0] _T_2891 = _T_2890 + _GEN_673; // @[PALU.scala 428:38]
  wire [6:0] _GEN_674 = {{6'd0}, _T_2869}; // @[PALU.scala 428:38]
  wire [7:0] _T_2892 = _T_2891 + _GEN_674; // @[PALU.scala 428:38]
  wire [7:0] _GEN_675 = {{7'd0}, _T_2871}; // @[PALU.scala 428:38]
  wire [8:0] _T_2893 = _T_2892 + _GEN_675; // @[PALU.scala 428:38]
  wire [8:0] _GEN_676 = {{8'd0}, _T_2873}; // @[PALU.scala 428:38]
  wire [9:0] _T_2894 = _T_2893 + _GEN_676; // @[PALU.scala 428:38]
  wire [9:0] _GEN_677 = {{9'd0}, _T_2875}; // @[PALU.scala 428:38]
  wire [10:0] _T_2895 = _T_2894 + _GEN_677; // @[PALU.scala 428:38]
  wire [10:0] _GEN_678 = {{10'd0}, _T_2877}; // @[PALU.scala 428:38]
  wire [11:0] _T_2896 = _T_2895 + _GEN_678; // @[PALU.scala 428:38]
  wire [11:0] _GEN_679 = {{11'd0}, _T_2879}; // @[PALU.scala 428:38]
  wire [12:0] _T_2897 = _T_2896 + _GEN_679; // @[PALU.scala 428:38]
  wire [12:0] _GEN_680 = {{12'd0}, _T_2881}; // @[PALU.scala 428:38]
  wire [13:0] _T_2898 = _T_2897 + _GEN_680; // @[PALU.scala 428:38]
  wire [13:0] _GEN_681 = {{13'd0}, _T_2883}; // @[PALU.scala 428:38]
  wire [14:0] _T_2899 = _T_2898 + _GEN_681; // @[PALU.scala 428:38]
  wire [14:0] _GEN_682 = {{14'd0}, _T_2885}; // @[PALU.scala 428:38]
  wire [15:0] _T_2900 = _T_2899 + _GEN_682; // @[PALU.scala 428:38]
  wire [15:0] _T_2902 = _T_2900 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_2903 = io_in_bits_DecodeIn_data_src2[0] ? _T_2900 : _T_2902; // @[PALU.scala 429:26]
  wire  _T_2906 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[47]; // @[PALU.scala 423:29]
  wire  _T_2908 = io_in_bits_DecodeIn_data_src1[32] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2910 = io_in_bits_DecodeIn_data_src1[33] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2912 = io_in_bits_DecodeIn_data_src1[34] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2914 = io_in_bits_DecodeIn_data_src1[35] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2916 = io_in_bits_DecodeIn_data_src1[36] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2918 = io_in_bits_DecodeIn_data_src1[37] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2920 = io_in_bits_DecodeIn_data_src1[38] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2922 = io_in_bits_DecodeIn_data_src1[39] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2924 = io_in_bits_DecodeIn_data_src1[40] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2926 = io_in_bits_DecodeIn_data_src1[41] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2928 = io_in_bits_DecodeIn_data_src1[42] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2930 = io_in_bits_DecodeIn_data_src1[43] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2932 = io_in_bits_DecodeIn_data_src1[44] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2934 = io_in_bits_DecodeIn_data_src1[45] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2936 = io_in_bits_DecodeIn_data_src1[46] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2938 = io_in_bits_DecodeIn_data_src1[47] == _T_2906; // @[PALU.scala 425:59]
  wire  _T_2940 = _T_2936 & _T_2938; // @[PALU.scala 427:113]
  wire  _T_2942 = _T_2934 & (_T_2936 & _T_2938); // @[PALU.scala 427:113]
  wire  _T_2944 = _T_2932 & (_T_2934 & (_T_2936 & _T_2938)); // @[PALU.scala 427:113]
  wire  _T_2946 = _T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))); // @[PALU.scala 427:113]
  wire  _T_2948 = _T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))); // @[PALU.scala 427:113]
  wire  _T_2950 = _T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))))); // @[PALU.scala 427:113]
  wire  _T_2952 = _T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))))); // @[PALU.scala 427:113]
  wire  _T_2954 = _T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))))))); // @[PALU.scala 427:113]
  wire  _T_2956 = _T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 &
    _T_2938)))))))); // @[PALU.scala 427:113]
  wire  _T_2958 = _T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (
    _T_2936 & _T_2938))))))))); // @[PALU.scala 427:113]
  wire  _T_2960 = _T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (
    _T_2934 & (_T_2936 & _T_2938)))))))))); // @[PALU.scala 427:113]
  wire  _T_2962 = _T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (_T_2930 & (
    _T_2932 & (_T_2934 & (_T_2936 & _T_2938))))))))))); // @[PALU.scala 427:113]
  wire  _T_2964 = _T_2912 & (_T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (_T_2928 & (
    _T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))))))))))); // @[PALU.scala 427:113]
  wire  _T_2966 = _T_2910 & (_T_2912 & (_T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (_T_2926 & (
    _T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938))))))))))))); // @[PALU.scala 427:113]
  wire  _T_2968 = _T_2908 & (_T_2910 & (_T_2912 & (_T_2914 & (_T_2916 & (_T_2918 & (_T_2920 & (_T_2922 & (_T_2924 & (
    _T_2926 & (_T_2928 & (_T_2930 & (_T_2932 & (_T_2934 & (_T_2936 & _T_2938)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_2969 = _T_2938 + _T_2940; // @[PALU.scala 428:38]
  wire [1:0] _GEN_683 = {{1'd0}, _T_2942}; // @[PALU.scala 428:38]
  wire [2:0] _T_2970 = _T_2969 + _GEN_683; // @[PALU.scala 428:38]
  wire [2:0] _GEN_684 = {{2'd0}, _T_2944}; // @[PALU.scala 428:38]
  wire [3:0] _T_2971 = _T_2970 + _GEN_684; // @[PALU.scala 428:38]
  wire [3:0] _GEN_685 = {{3'd0}, _T_2946}; // @[PALU.scala 428:38]
  wire [4:0] _T_2972 = _T_2971 + _GEN_685; // @[PALU.scala 428:38]
  wire [4:0] _GEN_686 = {{4'd0}, _T_2948}; // @[PALU.scala 428:38]
  wire [5:0] _T_2973 = _T_2972 + _GEN_686; // @[PALU.scala 428:38]
  wire [5:0] _GEN_687 = {{5'd0}, _T_2950}; // @[PALU.scala 428:38]
  wire [6:0] _T_2974 = _T_2973 + _GEN_687; // @[PALU.scala 428:38]
  wire [6:0] _GEN_688 = {{6'd0}, _T_2952}; // @[PALU.scala 428:38]
  wire [7:0] _T_2975 = _T_2974 + _GEN_688; // @[PALU.scala 428:38]
  wire [7:0] _GEN_689 = {{7'd0}, _T_2954}; // @[PALU.scala 428:38]
  wire [8:0] _T_2976 = _T_2975 + _GEN_689; // @[PALU.scala 428:38]
  wire [8:0] _GEN_690 = {{8'd0}, _T_2956}; // @[PALU.scala 428:38]
  wire [9:0] _T_2977 = _T_2976 + _GEN_690; // @[PALU.scala 428:38]
  wire [9:0] _GEN_691 = {{9'd0}, _T_2958}; // @[PALU.scala 428:38]
  wire [10:0] _T_2978 = _T_2977 + _GEN_691; // @[PALU.scala 428:38]
  wire [10:0] _GEN_692 = {{10'd0}, _T_2960}; // @[PALU.scala 428:38]
  wire [11:0] _T_2979 = _T_2978 + _GEN_692; // @[PALU.scala 428:38]
  wire [11:0] _GEN_693 = {{11'd0}, _T_2962}; // @[PALU.scala 428:38]
  wire [12:0] _T_2980 = _T_2979 + _GEN_693; // @[PALU.scala 428:38]
  wire [12:0] _GEN_694 = {{12'd0}, _T_2964}; // @[PALU.scala 428:38]
  wire [13:0] _T_2981 = _T_2980 + _GEN_694; // @[PALU.scala 428:38]
  wire [13:0] _GEN_695 = {{13'd0}, _T_2966}; // @[PALU.scala 428:38]
  wire [14:0] _T_2982 = _T_2981 + _GEN_695; // @[PALU.scala 428:38]
  wire [14:0] _GEN_696 = {{14'd0}, _T_2968}; // @[PALU.scala 428:38]
  wire [15:0] _T_2983 = _T_2982 + _GEN_696; // @[PALU.scala 428:38]
  wire [15:0] _T_2985 = _T_2983 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_2986 = io_in_bits_DecodeIn_data_src2[0] ? _T_2983 : _T_2985; // @[PALU.scala 429:26]
  wire  _T_2989 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[63]; // @[PALU.scala 423:29]
  wire  _T_2991 = io_in_bits_DecodeIn_data_src1[48] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2993 = io_in_bits_DecodeIn_data_src1[49] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2995 = io_in_bits_DecodeIn_data_src1[50] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2997 = io_in_bits_DecodeIn_data_src1[51] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_2999 = io_in_bits_DecodeIn_data_src1[52] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3001 = io_in_bits_DecodeIn_data_src1[53] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3003 = io_in_bits_DecodeIn_data_src1[54] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3005 = io_in_bits_DecodeIn_data_src1[55] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3007 = io_in_bits_DecodeIn_data_src1[56] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3009 = io_in_bits_DecodeIn_data_src1[57] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3011 = io_in_bits_DecodeIn_data_src1[58] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3013 = io_in_bits_DecodeIn_data_src1[59] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3015 = io_in_bits_DecodeIn_data_src1[60] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3017 = io_in_bits_DecodeIn_data_src1[61] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3019 = io_in_bits_DecodeIn_data_src1[62] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3021 = io_in_bits_DecodeIn_data_src1[63] == _T_2989; // @[PALU.scala 425:59]
  wire  _T_3023 = _T_3019 & _T_3021; // @[PALU.scala 427:113]
  wire  _T_3025 = _T_3017 & (_T_3019 & _T_3021); // @[PALU.scala 427:113]
  wire  _T_3027 = _T_3015 & (_T_3017 & (_T_3019 & _T_3021)); // @[PALU.scala 427:113]
  wire  _T_3029 = _T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))); // @[PALU.scala 427:113]
  wire  _T_3031 = _T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))); // @[PALU.scala 427:113]
  wire  _T_3033 = _T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))))); // @[PALU.scala 427:113]
  wire  _T_3035 = _T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))))); // @[PALU.scala 427:113]
  wire  _T_3037 = _T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))))))); // @[PALU.scala 427:113]
  wire  _T_3039 = _T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 &
    _T_3021)))))))); // @[PALU.scala 427:113]
  wire  _T_3041 = _T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (
    _T_3019 & _T_3021))))))))); // @[PALU.scala 427:113]
  wire  _T_3043 = _T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (
    _T_3017 & (_T_3019 & _T_3021)))))))))); // @[PALU.scala 427:113]
  wire  _T_3045 = _T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (_T_3013 & (
    _T_3015 & (_T_3017 & (_T_3019 & _T_3021))))))))))); // @[PALU.scala 427:113]
  wire  _T_3047 = _T_2995 & (_T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (_T_3011 & (
    _T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))))))))))); // @[PALU.scala 427:113]
  wire  _T_3049 = _T_2993 & (_T_2995 & (_T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (_T_3009 & (
    _T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3051 = _T_2991 & (_T_2993 & (_T_2995 & (_T_2997 & (_T_2999 & (_T_3001 & (_T_3003 & (_T_3005 & (_T_3007 & (
    _T_3009 & (_T_3011 & (_T_3013 & (_T_3015 & (_T_3017 & (_T_3019 & _T_3021)))))))))))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3052 = _T_3021 + _T_3023; // @[PALU.scala 428:38]
  wire [1:0] _GEN_697 = {{1'd0}, _T_3025}; // @[PALU.scala 428:38]
  wire [2:0] _T_3053 = _T_3052 + _GEN_697; // @[PALU.scala 428:38]
  wire [2:0] _GEN_698 = {{2'd0}, _T_3027}; // @[PALU.scala 428:38]
  wire [3:0] _T_3054 = _T_3053 + _GEN_698; // @[PALU.scala 428:38]
  wire [3:0] _GEN_699 = {{3'd0}, _T_3029}; // @[PALU.scala 428:38]
  wire [4:0] _T_3055 = _T_3054 + _GEN_699; // @[PALU.scala 428:38]
  wire [4:0] _GEN_700 = {{4'd0}, _T_3031}; // @[PALU.scala 428:38]
  wire [5:0] _T_3056 = _T_3055 + _GEN_700; // @[PALU.scala 428:38]
  wire [5:0] _GEN_701 = {{5'd0}, _T_3033}; // @[PALU.scala 428:38]
  wire [6:0] _T_3057 = _T_3056 + _GEN_701; // @[PALU.scala 428:38]
  wire [6:0] _GEN_702 = {{6'd0}, _T_3035}; // @[PALU.scala 428:38]
  wire [7:0] _T_3058 = _T_3057 + _GEN_702; // @[PALU.scala 428:38]
  wire [7:0] _GEN_703 = {{7'd0}, _T_3037}; // @[PALU.scala 428:38]
  wire [8:0] _T_3059 = _T_3058 + _GEN_703; // @[PALU.scala 428:38]
  wire [8:0] _GEN_704 = {{8'd0}, _T_3039}; // @[PALU.scala 428:38]
  wire [9:0] _T_3060 = _T_3059 + _GEN_704; // @[PALU.scala 428:38]
  wire [9:0] _GEN_705 = {{9'd0}, _T_3041}; // @[PALU.scala 428:38]
  wire [10:0] _T_3061 = _T_3060 + _GEN_705; // @[PALU.scala 428:38]
  wire [10:0] _GEN_706 = {{10'd0}, _T_3043}; // @[PALU.scala 428:38]
  wire [11:0] _T_3062 = _T_3061 + _GEN_706; // @[PALU.scala 428:38]
  wire [11:0] _GEN_707 = {{11'd0}, _T_3045}; // @[PALU.scala 428:38]
  wire [12:0] _T_3063 = _T_3062 + _GEN_707; // @[PALU.scala 428:38]
  wire [12:0] _GEN_708 = {{12'd0}, _T_3047}; // @[PALU.scala 428:38]
  wire [13:0] _T_3064 = _T_3063 + _GEN_708; // @[PALU.scala 428:38]
  wire [13:0] _GEN_709 = {{13'd0}, _T_3049}; // @[PALU.scala 428:38]
  wire [14:0] _T_3065 = _T_3064 + _GEN_709; // @[PALU.scala 428:38]
  wire [14:0] _GEN_710 = {{14'd0}, _T_3051}; // @[PALU.scala 428:38]
  wire [15:0] _T_3066 = _T_3065 + _GEN_710; // @[PALU.scala 428:38]
  wire [15:0] _T_3068 = _T_3066 - 16'h1; // @[PALU.scala 429:44]
  wire [15:0] _T_3069 = io_in_bits_DecodeIn_data_src2[0] ? _T_3066 : _T_3068; // @[PALU.scala 429:26]
  wire [63:0] _T_3072 = {_T_3069,_T_2986,_T_2903,_T_2820}; // @[Cat.scala 30:58]
  wire  _T_3077 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[7]; // @[PALU.scala 423:29]
  wire  _T_3079 = io_in_bits_DecodeIn_data_src1[0] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3081 = io_in_bits_DecodeIn_data_src1[1] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3083 = io_in_bits_DecodeIn_data_src1[2] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3085 = io_in_bits_DecodeIn_data_src1[3] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3087 = io_in_bits_DecodeIn_data_src1[4] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3089 = io_in_bits_DecodeIn_data_src1[5] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3091 = io_in_bits_DecodeIn_data_src1[6] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3093 = io_in_bits_DecodeIn_data_src1[7] == _T_3077; // @[PALU.scala 425:59]
  wire  _T_3095 = _T_3091 & _T_3093; // @[PALU.scala 427:113]
  wire  _T_3097 = _T_3089 & (_T_3091 & _T_3093); // @[PALU.scala 427:113]
  wire  _T_3099 = _T_3087 & (_T_3089 & (_T_3091 & _T_3093)); // @[PALU.scala 427:113]
  wire  _T_3101 = _T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093))); // @[PALU.scala 427:113]
  wire  _T_3103 = _T_3083 & (_T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093)))); // @[PALU.scala 427:113]
  wire  _T_3105 = _T_3081 & (_T_3083 & (_T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093))))); // @[PALU.scala 427:113]
  wire  _T_3107 = _T_3079 & (_T_3081 & (_T_3083 & (_T_3085 & (_T_3087 & (_T_3089 & (_T_3091 & _T_3093)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3108 = _T_3093 + _T_3095; // @[PALU.scala 428:38]
  wire [1:0] _GEN_711 = {{1'd0}, _T_3097}; // @[PALU.scala 428:38]
  wire [2:0] _T_3109 = _T_3108 + _GEN_711; // @[PALU.scala 428:38]
  wire [2:0] _GEN_712 = {{2'd0}, _T_3099}; // @[PALU.scala 428:38]
  wire [3:0] _T_3110 = _T_3109 + _GEN_712; // @[PALU.scala 428:38]
  wire [3:0] _GEN_713 = {{3'd0}, _T_3101}; // @[PALU.scala 428:38]
  wire [4:0] _T_3111 = _T_3110 + _GEN_713; // @[PALU.scala 428:38]
  wire [4:0] _GEN_714 = {{4'd0}, _T_3103}; // @[PALU.scala 428:38]
  wire [5:0] _T_3112 = _T_3111 + _GEN_714; // @[PALU.scala 428:38]
  wire [5:0] _GEN_715 = {{5'd0}, _T_3105}; // @[PALU.scala 428:38]
  wire [6:0] _T_3113 = _T_3112 + _GEN_715; // @[PALU.scala 428:38]
  wire [6:0] _GEN_716 = {{6'd0}, _T_3107}; // @[PALU.scala 428:38]
  wire [7:0] _T_3114 = _T_3113 + _GEN_716; // @[PALU.scala 428:38]
  wire [7:0] _T_3116 = _T_3114 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3117 = io_in_bits_DecodeIn_data_src2[0] ? _T_3114 : _T_3116; // @[PALU.scala 429:26]
  wire  _T_3120 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[15]; // @[PALU.scala 423:29]
  wire  _T_3122 = io_in_bits_DecodeIn_data_src1[8] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3124 = io_in_bits_DecodeIn_data_src1[9] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3126 = io_in_bits_DecodeIn_data_src1[10] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3128 = io_in_bits_DecodeIn_data_src1[11] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3130 = io_in_bits_DecodeIn_data_src1[12] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3132 = io_in_bits_DecodeIn_data_src1[13] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3134 = io_in_bits_DecodeIn_data_src1[14] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3136 = io_in_bits_DecodeIn_data_src1[15] == _T_3120; // @[PALU.scala 425:59]
  wire  _T_3138 = _T_3134 & _T_3136; // @[PALU.scala 427:113]
  wire  _T_3140 = _T_3132 & (_T_3134 & _T_3136); // @[PALU.scala 427:113]
  wire  _T_3142 = _T_3130 & (_T_3132 & (_T_3134 & _T_3136)); // @[PALU.scala 427:113]
  wire  _T_3144 = _T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136))); // @[PALU.scala 427:113]
  wire  _T_3146 = _T_3126 & (_T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136)))); // @[PALU.scala 427:113]
  wire  _T_3148 = _T_3124 & (_T_3126 & (_T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136))))); // @[PALU.scala 427:113]
  wire  _T_3150 = _T_3122 & (_T_3124 & (_T_3126 & (_T_3128 & (_T_3130 & (_T_3132 & (_T_3134 & _T_3136)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3151 = _T_3136 + _T_3138; // @[PALU.scala 428:38]
  wire [1:0] _GEN_717 = {{1'd0}, _T_3140}; // @[PALU.scala 428:38]
  wire [2:0] _T_3152 = _T_3151 + _GEN_717; // @[PALU.scala 428:38]
  wire [2:0] _GEN_718 = {{2'd0}, _T_3142}; // @[PALU.scala 428:38]
  wire [3:0] _T_3153 = _T_3152 + _GEN_718; // @[PALU.scala 428:38]
  wire [3:0] _GEN_719 = {{3'd0}, _T_3144}; // @[PALU.scala 428:38]
  wire [4:0] _T_3154 = _T_3153 + _GEN_719; // @[PALU.scala 428:38]
  wire [4:0] _GEN_720 = {{4'd0}, _T_3146}; // @[PALU.scala 428:38]
  wire [5:0] _T_3155 = _T_3154 + _GEN_720; // @[PALU.scala 428:38]
  wire [5:0] _GEN_721 = {{5'd0}, _T_3148}; // @[PALU.scala 428:38]
  wire [6:0] _T_3156 = _T_3155 + _GEN_721; // @[PALU.scala 428:38]
  wire [6:0] _GEN_722 = {{6'd0}, _T_3150}; // @[PALU.scala 428:38]
  wire [7:0] _T_3157 = _T_3156 + _GEN_722; // @[PALU.scala 428:38]
  wire [7:0] _T_3159 = _T_3157 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3160 = io_in_bits_DecodeIn_data_src2[0] ? _T_3157 : _T_3159; // @[PALU.scala 429:26]
  wire  _T_3163 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[23]; // @[PALU.scala 423:29]
  wire  _T_3165 = io_in_bits_DecodeIn_data_src1[16] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3167 = io_in_bits_DecodeIn_data_src1[17] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3169 = io_in_bits_DecodeIn_data_src1[18] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3171 = io_in_bits_DecodeIn_data_src1[19] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3173 = io_in_bits_DecodeIn_data_src1[20] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3175 = io_in_bits_DecodeIn_data_src1[21] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3177 = io_in_bits_DecodeIn_data_src1[22] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3179 = io_in_bits_DecodeIn_data_src1[23] == _T_3163; // @[PALU.scala 425:59]
  wire  _T_3181 = _T_3177 & _T_3179; // @[PALU.scala 427:113]
  wire  _T_3183 = _T_3175 & (_T_3177 & _T_3179); // @[PALU.scala 427:113]
  wire  _T_3185 = _T_3173 & (_T_3175 & (_T_3177 & _T_3179)); // @[PALU.scala 427:113]
  wire  _T_3187 = _T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179))); // @[PALU.scala 427:113]
  wire  _T_3189 = _T_3169 & (_T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179)))); // @[PALU.scala 427:113]
  wire  _T_3191 = _T_3167 & (_T_3169 & (_T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179))))); // @[PALU.scala 427:113]
  wire  _T_3193 = _T_3165 & (_T_3167 & (_T_3169 & (_T_3171 & (_T_3173 & (_T_3175 & (_T_3177 & _T_3179)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3194 = _T_3179 + _T_3181; // @[PALU.scala 428:38]
  wire [1:0] _GEN_723 = {{1'd0}, _T_3183}; // @[PALU.scala 428:38]
  wire [2:0] _T_3195 = _T_3194 + _GEN_723; // @[PALU.scala 428:38]
  wire [2:0] _GEN_724 = {{2'd0}, _T_3185}; // @[PALU.scala 428:38]
  wire [3:0] _T_3196 = _T_3195 + _GEN_724; // @[PALU.scala 428:38]
  wire [3:0] _GEN_725 = {{3'd0}, _T_3187}; // @[PALU.scala 428:38]
  wire [4:0] _T_3197 = _T_3196 + _GEN_725; // @[PALU.scala 428:38]
  wire [4:0] _GEN_726 = {{4'd0}, _T_3189}; // @[PALU.scala 428:38]
  wire [5:0] _T_3198 = _T_3197 + _GEN_726; // @[PALU.scala 428:38]
  wire [5:0] _GEN_727 = {{5'd0}, _T_3191}; // @[PALU.scala 428:38]
  wire [6:0] _T_3199 = _T_3198 + _GEN_727; // @[PALU.scala 428:38]
  wire [6:0] _GEN_728 = {{6'd0}, _T_3193}; // @[PALU.scala 428:38]
  wire [7:0] _T_3200 = _T_3199 + _GEN_728; // @[PALU.scala 428:38]
  wire [7:0] _T_3202 = _T_3200 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3203 = io_in_bits_DecodeIn_data_src2[0] ? _T_3200 : _T_3202; // @[PALU.scala 429:26]
  wire  _T_3206 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[31]; // @[PALU.scala 423:29]
  wire  _T_3208 = io_in_bits_DecodeIn_data_src1[24] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3210 = io_in_bits_DecodeIn_data_src1[25] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3212 = io_in_bits_DecodeIn_data_src1[26] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3214 = io_in_bits_DecodeIn_data_src1[27] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3216 = io_in_bits_DecodeIn_data_src1[28] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3218 = io_in_bits_DecodeIn_data_src1[29] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3220 = io_in_bits_DecodeIn_data_src1[30] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3222 = io_in_bits_DecodeIn_data_src1[31] == _T_3206; // @[PALU.scala 425:59]
  wire  _T_3224 = _T_3220 & _T_3222; // @[PALU.scala 427:113]
  wire  _T_3226 = _T_3218 & (_T_3220 & _T_3222); // @[PALU.scala 427:113]
  wire  _T_3228 = _T_3216 & (_T_3218 & (_T_3220 & _T_3222)); // @[PALU.scala 427:113]
  wire  _T_3230 = _T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222))); // @[PALU.scala 427:113]
  wire  _T_3232 = _T_3212 & (_T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222)))); // @[PALU.scala 427:113]
  wire  _T_3234 = _T_3210 & (_T_3212 & (_T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222))))); // @[PALU.scala 427:113]
  wire  _T_3236 = _T_3208 & (_T_3210 & (_T_3212 & (_T_3214 & (_T_3216 & (_T_3218 & (_T_3220 & _T_3222)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3237 = _T_3222 + _T_3224; // @[PALU.scala 428:38]
  wire [1:0] _GEN_729 = {{1'd0}, _T_3226}; // @[PALU.scala 428:38]
  wire [2:0] _T_3238 = _T_3237 + _GEN_729; // @[PALU.scala 428:38]
  wire [2:0] _GEN_730 = {{2'd0}, _T_3228}; // @[PALU.scala 428:38]
  wire [3:0] _T_3239 = _T_3238 + _GEN_730; // @[PALU.scala 428:38]
  wire [3:0] _GEN_731 = {{3'd0}, _T_3230}; // @[PALU.scala 428:38]
  wire [4:0] _T_3240 = _T_3239 + _GEN_731; // @[PALU.scala 428:38]
  wire [4:0] _GEN_732 = {{4'd0}, _T_3232}; // @[PALU.scala 428:38]
  wire [5:0] _T_3241 = _T_3240 + _GEN_732; // @[PALU.scala 428:38]
  wire [5:0] _GEN_733 = {{5'd0}, _T_3234}; // @[PALU.scala 428:38]
  wire [6:0] _T_3242 = _T_3241 + _GEN_733; // @[PALU.scala 428:38]
  wire [6:0] _GEN_734 = {{6'd0}, _T_3236}; // @[PALU.scala 428:38]
  wire [7:0] _T_3243 = _T_3242 + _GEN_734; // @[PALU.scala 428:38]
  wire [7:0] _T_3245 = _T_3243 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3246 = io_in_bits_DecodeIn_data_src2[0] ? _T_3243 : _T_3245; // @[PALU.scala 429:26]
  wire  _T_3249 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[39]; // @[PALU.scala 423:29]
  wire  _T_3251 = io_in_bits_DecodeIn_data_src1[32] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3253 = io_in_bits_DecodeIn_data_src1[33] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3255 = io_in_bits_DecodeIn_data_src1[34] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3257 = io_in_bits_DecodeIn_data_src1[35] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3259 = io_in_bits_DecodeIn_data_src1[36] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3261 = io_in_bits_DecodeIn_data_src1[37] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3263 = io_in_bits_DecodeIn_data_src1[38] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3265 = io_in_bits_DecodeIn_data_src1[39] == _T_3249; // @[PALU.scala 425:59]
  wire  _T_3267 = _T_3263 & _T_3265; // @[PALU.scala 427:113]
  wire  _T_3269 = _T_3261 & (_T_3263 & _T_3265); // @[PALU.scala 427:113]
  wire  _T_3271 = _T_3259 & (_T_3261 & (_T_3263 & _T_3265)); // @[PALU.scala 427:113]
  wire  _T_3273 = _T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265))); // @[PALU.scala 427:113]
  wire  _T_3275 = _T_3255 & (_T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265)))); // @[PALU.scala 427:113]
  wire  _T_3277 = _T_3253 & (_T_3255 & (_T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265))))); // @[PALU.scala 427:113]
  wire  _T_3279 = _T_3251 & (_T_3253 & (_T_3255 & (_T_3257 & (_T_3259 & (_T_3261 & (_T_3263 & _T_3265)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3280 = _T_3265 + _T_3267; // @[PALU.scala 428:38]
  wire [1:0] _GEN_735 = {{1'd0}, _T_3269}; // @[PALU.scala 428:38]
  wire [2:0] _T_3281 = _T_3280 + _GEN_735; // @[PALU.scala 428:38]
  wire [2:0] _GEN_736 = {{2'd0}, _T_3271}; // @[PALU.scala 428:38]
  wire [3:0] _T_3282 = _T_3281 + _GEN_736; // @[PALU.scala 428:38]
  wire [3:0] _GEN_737 = {{3'd0}, _T_3273}; // @[PALU.scala 428:38]
  wire [4:0] _T_3283 = _T_3282 + _GEN_737; // @[PALU.scala 428:38]
  wire [4:0] _GEN_738 = {{4'd0}, _T_3275}; // @[PALU.scala 428:38]
  wire [5:0] _T_3284 = _T_3283 + _GEN_738; // @[PALU.scala 428:38]
  wire [5:0] _GEN_739 = {{5'd0}, _T_3277}; // @[PALU.scala 428:38]
  wire [6:0] _T_3285 = _T_3284 + _GEN_739; // @[PALU.scala 428:38]
  wire [6:0] _GEN_740 = {{6'd0}, _T_3279}; // @[PALU.scala 428:38]
  wire [7:0] _T_3286 = _T_3285 + _GEN_740; // @[PALU.scala 428:38]
  wire [7:0] _T_3288 = _T_3286 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3289 = io_in_bits_DecodeIn_data_src2[0] ? _T_3286 : _T_3288; // @[PALU.scala 429:26]
  wire  _T_3292 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[47]; // @[PALU.scala 423:29]
  wire  _T_3294 = io_in_bits_DecodeIn_data_src1[40] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3296 = io_in_bits_DecodeIn_data_src1[41] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3298 = io_in_bits_DecodeIn_data_src1[42] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3300 = io_in_bits_DecodeIn_data_src1[43] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3302 = io_in_bits_DecodeIn_data_src1[44] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3304 = io_in_bits_DecodeIn_data_src1[45] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3306 = io_in_bits_DecodeIn_data_src1[46] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3308 = io_in_bits_DecodeIn_data_src1[47] == _T_3292; // @[PALU.scala 425:59]
  wire  _T_3310 = _T_3306 & _T_3308; // @[PALU.scala 427:113]
  wire  _T_3312 = _T_3304 & (_T_3306 & _T_3308); // @[PALU.scala 427:113]
  wire  _T_3314 = _T_3302 & (_T_3304 & (_T_3306 & _T_3308)); // @[PALU.scala 427:113]
  wire  _T_3316 = _T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308))); // @[PALU.scala 427:113]
  wire  _T_3318 = _T_3298 & (_T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308)))); // @[PALU.scala 427:113]
  wire  _T_3320 = _T_3296 & (_T_3298 & (_T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308))))); // @[PALU.scala 427:113]
  wire  _T_3322 = _T_3294 & (_T_3296 & (_T_3298 & (_T_3300 & (_T_3302 & (_T_3304 & (_T_3306 & _T_3308)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3323 = _T_3308 + _T_3310; // @[PALU.scala 428:38]
  wire [1:0] _GEN_741 = {{1'd0}, _T_3312}; // @[PALU.scala 428:38]
  wire [2:0] _T_3324 = _T_3323 + _GEN_741; // @[PALU.scala 428:38]
  wire [2:0] _GEN_742 = {{2'd0}, _T_3314}; // @[PALU.scala 428:38]
  wire [3:0] _T_3325 = _T_3324 + _GEN_742; // @[PALU.scala 428:38]
  wire [3:0] _GEN_743 = {{3'd0}, _T_3316}; // @[PALU.scala 428:38]
  wire [4:0] _T_3326 = _T_3325 + _GEN_743; // @[PALU.scala 428:38]
  wire [4:0] _GEN_744 = {{4'd0}, _T_3318}; // @[PALU.scala 428:38]
  wire [5:0] _T_3327 = _T_3326 + _GEN_744; // @[PALU.scala 428:38]
  wire [5:0] _GEN_745 = {{5'd0}, _T_3320}; // @[PALU.scala 428:38]
  wire [6:0] _T_3328 = _T_3327 + _GEN_745; // @[PALU.scala 428:38]
  wire [6:0] _GEN_746 = {{6'd0}, _T_3322}; // @[PALU.scala 428:38]
  wire [7:0] _T_3329 = _T_3328 + _GEN_746; // @[PALU.scala 428:38]
  wire [7:0] _T_3331 = _T_3329 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3332 = io_in_bits_DecodeIn_data_src2[0] ? _T_3329 : _T_3331; // @[PALU.scala 429:26]
  wire  _T_3335 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[55]; // @[PALU.scala 423:29]
  wire  _T_3337 = io_in_bits_DecodeIn_data_src1[48] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3339 = io_in_bits_DecodeIn_data_src1[49] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3341 = io_in_bits_DecodeIn_data_src1[50] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3343 = io_in_bits_DecodeIn_data_src1[51] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3345 = io_in_bits_DecodeIn_data_src1[52] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3347 = io_in_bits_DecodeIn_data_src1[53] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3349 = io_in_bits_DecodeIn_data_src1[54] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3351 = io_in_bits_DecodeIn_data_src1[55] == _T_3335; // @[PALU.scala 425:59]
  wire  _T_3353 = _T_3349 & _T_3351; // @[PALU.scala 427:113]
  wire  _T_3355 = _T_3347 & (_T_3349 & _T_3351); // @[PALU.scala 427:113]
  wire  _T_3357 = _T_3345 & (_T_3347 & (_T_3349 & _T_3351)); // @[PALU.scala 427:113]
  wire  _T_3359 = _T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351))); // @[PALU.scala 427:113]
  wire  _T_3361 = _T_3341 & (_T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351)))); // @[PALU.scala 427:113]
  wire  _T_3363 = _T_3339 & (_T_3341 & (_T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351))))); // @[PALU.scala 427:113]
  wire  _T_3365 = _T_3337 & (_T_3339 & (_T_3341 & (_T_3343 & (_T_3345 & (_T_3347 & (_T_3349 & _T_3351)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3366 = _T_3351 + _T_3353; // @[PALU.scala 428:38]
  wire [1:0] _GEN_747 = {{1'd0}, _T_3355}; // @[PALU.scala 428:38]
  wire [2:0] _T_3367 = _T_3366 + _GEN_747; // @[PALU.scala 428:38]
  wire [2:0] _GEN_748 = {{2'd0}, _T_3357}; // @[PALU.scala 428:38]
  wire [3:0] _T_3368 = _T_3367 + _GEN_748; // @[PALU.scala 428:38]
  wire [3:0] _GEN_749 = {{3'd0}, _T_3359}; // @[PALU.scala 428:38]
  wire [4:0] _T_3369 = _T_3368 + _GEN_749; // @[PALU.scala 428:38]
  wire [4:0] _GEN_750 = {{4'd0}, _T_3361}; // @[PALU.scala 428:38]
  wire [5:0] _T_3370 = _T_3369 + _GEN_750; // @[PALU.scala 428:38]
  wire [5:0] _GEN_751 = {{5'd0}, _T_3363}; // @[PALU.scala 428:38]
  wire [6:0] _T_3371 = _T_3370 + _GEN_751; // @[PALU.scala 428:38]
  wire [6:0] _GEN_752 = {{6'd0}, _T_3365}; // @[PALU.scala 428:38]
  wire [7:0] _T_3372 = _T_3371 + _GEN_752; // @[PALU.scala 428:38]
  wire [7:0] _T_3374 = _T_3372 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3375 = io_in_bits_DecodeIn_data_src2[0] ? _T_3372 : _T_3374; // @[PALU.scala 429:26]
  wire  _T_3378 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[63]; // @[PALU.scala 423:29]
  wire  _T_3380 = io_in_bits_DecodeIn_data_src1[56] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3382 = io_in_bits_DecodeIn_data_src1[57] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3384 = io_in_bits_DecodeIn_data_src1[58] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3386 = io_in_bits_DecodeIn_data_src1[59] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3388 = io_in_bits_DecodeIn_data_src1[60] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3390 = io_in_bits_DecodeIn_data_src1[61] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3392 = io_in_bits_DecodeIn_data_src1[62] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3394 = io_in_bits_DecodeIn_data_src1[63] == _T_3378; // @[PALU.scala 425:59]
  wire  _T_3396 = _T_3392 & _T_3394; // @[PALU.scala 427:113]
  wire  _T_3398 = _T_3390 & (_T_3392 & _T_3394); // @[PALU.scala 427:113]
  wire  _T_3400 = _T_3388 & (_T_3390 & (_T_3392 & _T_3394)); // @[PALU.scala 427:113]
  wire  _T_3402 = _T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394))); // @[PALU.scala 427:113]
  wire  _T_3404 = _T_3384 & (_T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394)))); // @[PALU.scala 427:113]
  wire  _T_3406 = _T_3382 & (_T_3384 & (_T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394))))); // @[PALU.scala 427:113]
  wire  _T_3408 = _T_3380 & (_T_3382 & (_T_3384 & (_T_3386 & (_T_3388 & (_T_3390 & (_T_3392 & _T_3394)))))); // @[PALU.scala 427:113]
  wire [1:0] _T_3409 = _T_3394 + _T_3396; // @[PALU.scala 428:38]
  wire [1:0] _GEN_753 = {{1'd0}, _T_3398}; // @[PALU.scala 428:38]
  wire [2:0] _T_3410 = _T_3409 + _GEN_753; // @[PALU.scala 428:38]
  wire [2:0] _GEN_754 = {{2'd0}, _T_3400}; // @[PALU.scala 428:38]
  wire [3:0] _T_3411 = _T_3410 + _GEN_754; // @[PALU.scala 428:38]
  wire [3:0] _GEN_755 = {{3'd0}, _T_3402}; // @[PALU.scala 428:38]
  wire [4:0] _T_3412 = _T_3411 + _GEN_755; // @[PALU.scala 428:38]
  wire [4:0] _GEN_756 = {{4'd0}, _T_3404}; // @[PALU.scala 428:38]
  wire [5:0] _T_3413 = _T_3412 + _GEN_756; // @[PALU.scala 428:38]
  wire [5:0] _GEN_757 = {{5'd0}, _T_3406}; // @[PALU.scala 428:38]
  wire [6:0] _T_3414 = _T_3413 + _GEN_757; // @[PALU.scala 428:38]
  wire [6:0] _GEN_758 = {{6'd0}, _T_3408}; // @[PALU.scala 428:38]
  wire [7:0] _T_3415 = _T_3414 + _GEN_758; // @[PALU.scala 428:38]
  wire [7:0] _T_3417 = _T_3415 - 8'h1; // @[PALU.scala 429:44]
  wire [7:0] _T_3418 = io_in_bits_DecodeIn_data_src2[0] ? _T_3415 : _T_3417; // @[PALU.scala 429:26]
  wire [63:0] _T_3425 = {_T_3418,_T_3375,_T_3332,_T_3289,_T_3246,_T_3203,_T_3160,_T_3117}; // @[Cat.scala 30:58]
  wire  _T_3430 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[31]; // @[PALU.scala 423:29]
  wire  _T_3432 = io_in_bits_DecodeIn_data_src1[0] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3434 = io_in_bits_DecodeIn_data_src1[1] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3436 = io_in_bits_DecodeIn_data_src1[2] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3438 = io_in_bits_DecodeIn_data_src1[3] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3440 = io_in_bits_DecodeIn_data_src1[4] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3442 = io_in_bits_DecodeIn_data_src1[5] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3444 = io_in_bits_DecodeIn_data_src1[6] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3446 = io_in_bits_DecodeIn_data_src1[7] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3448 = io_in_bits_DecodeIn_data_src1[8] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3450 = io_in_bits_DecodeIn_data_src1[9] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3452 = io_in_bits_DecodeIn_data_src1[10] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3454 = io_in_bits_DecodeIn_data_src1[11] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3456 = io_in_bits_DecodeIn_data_src1[12] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3458 = io_in_bits_DecodeIn_data_src1[13] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3460 = io_in_bits_DecodeIn_data_src1[14] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3462 = io_in_bits_DecodeIn_data_src1[15] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3464 = io_in_bits_DecodeIn_data_src1[16] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3466 = io_in_bits_DecodeIn_data_src1[17] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3468 = io_in_bits_DecodeIn_data_src1[18] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3470 = io_in_bits_DecodeIn_data_src1[19] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3472 = io_in_bits_DecodeIn_data_src1[20] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3474 = io_in_bits_DecodeIn_data_src1[21] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3476 = io_in_bits_DecodeIn_data_src1[22] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3478 = io_in_bits_DecodeIn_data_src1[23] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3480 = io_in_bits_DecodeIn_data_src1[24] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3482 = io_in_bits_DecodeIn_data_src1[25] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3484 = io_in_bits_DecodeIn_data_src1[26] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3486 = io_in_bits_DecodeIn_data_src1[27] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3488 = io_in_bits_DecodeIn_data_src1[28] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3490 = io_in_bits_DecodeIn_data_src1[29] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3492 = io_in_bits_DecodeIn_data_src1[30] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3494 = io_in_bits_DecodeIn_data_src1[31] == _T_3430; // @[PALU.scala 425:59]
  wire  _T_3496 = _T_3492 & _T_3494; // @[PALU.scala 427:113]
  wire  _T_3498 = _T_3490 & (_T_3492 & _T_3494); // @[PALU.scala 427:113]
  wire  _T_3500 = _T_3488 & (_T_3490 & (_T_3492 & _T_3494)); // @[PALU.scala 427:113]
  wire  _T_3502 = _T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))); // @[PALU.scala 427:113]
  wire  _T_3504 = _T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))); // @[PALU.scala 427:113]
  wire  _T_3506 = _T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))); // @[PALU.scala 427:113]
  wire  _T_3508 = _T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))); // @[PALU.scala 427:113]
  wire  _T_3510 = _T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))); // @[PALU.scala 427:113]
  wire  _T_3512 = _T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 &
    _T_3494)))))))); // @[PALU.scala 427:113]
  wire  _T_3514 = _T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (
    _T_3492 & _T_3494))))))))); // @[PALU.scala 427:113]
  wire  _T_3516 = _T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (
    _T_3490 & (_T_3492 & _T_3494)))))))))); // @[PALU.scala 427:113]
  wire  _T_3518 = _T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (
    _T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))); // @[PALU.scala 427:113]
  wire  _T_3520 = _T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (
    _T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))); // @[PALU.scala 427:113]
  wire  _T_3522 = _T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (
    _T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3524 = _T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (
    _T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3526 = _T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (
    _T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3528 = _T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (
    _T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3530 = _T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (
    _T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))
    )))))); // @[PALU.scala 427:113]
  wire  _T_3532 = _T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (
    _T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494
    )))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3534 = _T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (
    _T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (
    _T_3492 & _T_3494))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3536 = _T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (
    _T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (
    _T_3490 & (_T_3492 & _T_3494)))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3538 = _T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (
    _T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (
    _T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3540 = _T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (
    _T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (
    _T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3542 = _T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (
    _T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (
    _T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3544 = _T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (
    _T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (
    _T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3546 = _T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (
    _T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (
    _T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3548 = _T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (_T_3456 & (
    _T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (_T_3476 & (
    _T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494))))))))))))))))))))))
    )))); // @[PALU.scala 427:113]
  wire  _T_3550 = _T_3438 & (_T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (_T_3454 & (
    _T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (_T_3474 & (
    _T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494)))))))))))
    )))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3552 = _T_3436 & (_T_3438 & (_T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (_T_3452 & (
    _T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (_T_3472 & (
    _T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (_T_3492 & _T_3494
    )))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3554 = _T_3434 & (_T_3436 & (_T_3438 & (_T_3440 & (_T_3442 & (_T_3444 & (_T_3446 & (_T_3448 & (_T_3450 & (
    _T_3452 & (_T_3454 & (_T_3456 & (_T_3458 & (_T_3460 & (_T_3462 & (_T_3464 & (_T_3466 & (_T_3468 & (_T_3470 & (
    _T_3472 & (_T_3474 & (_T_3476 & (_T_3478 & (_T_3480 & (_T_3482 & (_T_3484 & (_T_3486 & (_T_3488 & (_T_3490 & (
    _T_3492 & _T_3494))))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3556 = _T_3432 & _T_3554; // @[PALU.scala 427:113]
  wire [1:0] _T_3557 = _T_3494 + _T_3496; // @[PALU.scala 428:38]
  wire [1:0] _GEN_759 = {{1'd0}, _T_3498}; // @[PALU.scala 428:38]
  wire [2:0] _T_3558 = _T_3557 + _GEN_759; // @[PALU.scala 428:38]
  wire [2:0] _GEN_760 = {{2'd0}, _T_3500}; // @[PALU.scala 428:38]
  wire [3:0] _T_3559 = _T_3558 + _GEN_760; // @[PALU.scala 428:38]
  wire [3:0] _GEN_761 = {{3'd0}, _T_3502}; // @[PALU.scala 428:38]
  wire [4:0] _T_3560 = _T_3559 + _GEN_761; // @[PALU.scala 428:38]
  wire [4:0] _GEN_762 = {{4'd0}, _T_3504}; // @[PALU.scala 428:38]
  wire [5:0] _T_3561 = _T_3560 + _GEN_762; // @[PALU.scala 428:38]
  wire [5:0] _GEN_763 = {{5'd0}, _T_3506}; // @[PALU.scala 428:38]
  wire [6:0] _T_3562 = _T_3561 + _GEN_763; // @[PALU.scala 428:38]
  wire [6:0] _GEN_764 = {{6'd0}, _T_3508}; // @[PALU.scala 428:38]
  wire [7:0] _T_3563 = _T_3562 + _GEN_764; // @[PALU.scala 428:38]
  wire [7:0] _GEN_765 = {{7'd0}, _T_3510}; // @[PALU.scala 428:38]
  wire [8:0] _T_3564 = _T_3563 + _GEN_765; // @[PALU.scala 428:38]
  wire [8:0] _GEN_766 = {{8'd0}, _T_3512}; // @[PALU.scala 428:38]
  wire [9:0] _T_3565 = _T_3564 + _GEN_766; // @[PALU.scala 428:38]
  wire [9:0] _GEN_767 = {{9'd0}, _T_3514}; // @[PALU.scala 428:38]
  wire [10:0] _T_3566 = _T_3565 + _GEN_767; // @[PALU.scala 428:38]
  wire [10:0] _GEN_768 = {{10'd0}, _T_3516}; // @[PALU.scala 428:38]
  wire [11:0] _T_3567 = _T_3566 + _GEN_768; // @[PALU.scala 428:38]
  wire [11:0] _GEN_769 = {{11'd0}, _T_3518}; // @[PALU.scala 428:38]
  wire [12:0] _T_3568 = _T_3567 + _GEN_769; // @[PALU.scala 428:38]
  wire [12:0] _GEN_770 = {{12'd0}, _T_3520}; // @[PALU.scala 428:38]
  wire [13:0] _T_3569 = _T_3568 + _GEN_770; // @[PALU.scala 428:38]
  wire [13:0] _GEN_771 = {{13'd0}, _T_3522}; // @[PALU.scala 428:38]
  wire [14:0] _T_3570 = _T_3569 + _GEN_771; // @[PALU.scala 428:38]
  wire [14:0] _GEN_772 = {{14'd0}, _T_3524}; // @[PALU.scala 428:38]
  wire [15:0] _T_3571 = _T_3570 + _GEN_772; // @[PALU.scala 428:38]
  wire [15:0] _GEN_773 = {{15'd0}, _T_3526}; // @[PALU.scala 428:38]
  wire [16:0] _T_3572 = _T_3571 + _GEN_773; // @[PALU.scala 428:38]
  wire [16:0] _GEN_774 = {{16'd0}, _T_3528}; // @[PALU.scala 428:38]
  wire [17:0] _T_3573 = _T_3572 + _GEN_774; // @[PALU.scala 428:38]
  wire [17:0] _GEN_775 = {{17'd0}, _T_3530}; // @[PALU.scala 428:38]
  wire [18:0] _T_3574 = _T_3573 + _GEN_775; // @[PALU.scala 428:38]
  wire [18:0] _GEN_776 = {{18'd0}, _T_3532}; // @[PALU.scala 428:38]
  wire [19:0] _T_3575 = _T_3574 + _GEN_776; // @[PALU.scala 428:38]
  wire [19:0] _GEN_777 = {{19'd0}, _T_3534}; // @[PALU.scala 428:38]
  wire [20:0] _T_3576 = _T_3575 + _GEN_777; // @[PALU.scala 428:38]
  wire [20:0] _GEN_778 = {{20'd0}, _T_3536}; // @[PALU.scala 428:38]
  wire [21:0] _T_3577 = _T_3576 + _GEN_778; // @[PALU.scala 428:38]
  wire [21:0] _GEN_779 = {{21'd0}, _T_3538}; // @[PALU.scala 428:38]
  wire [22:0] _T_3578 = _T_3577 + _GEN_779; // @[PALU.scala 428:38]
  wire [22:0] _GEN_780 = {{22'd0}, _T_3540}; // @[PALU.scala 428:38]
  wire [23:0] _T_3579 = _T_3578 + _GEN_780; // @[PALU.scala 428:38]
  wire [23:0] _GEN_781 = {{23'd0}, _T_3542}; // @[PALU.scala 428:38]
  wire [24:0] _T_3580 = _T_3579 + _GEN_781; // @[PALU.scala 428:38]
  wire [24:0] _GEN_782 = {{24'd0}, _T_3544}; // @[PALU.scala 428:38]
  wire [25:0] _T_3581 = _T_3580 + _GEN_782; // @[PALU.scala 428:38]
  wire [25:0] _GEN_783 = {{25'd0}, _T_3546}; // @[PALU.scala 428:38]
  wire [26:0] _T_3582 = _T_3581 + _GEN_783; // @[PALU.scala 428:38]
  wire [26:0] _GEN_784 = {{26'd0}, _T_3548}; // @[PALU.scala 428:38]
  wire [27:0] _T_3583 = _T_3582 + _GEN_784; // @[PALU.scala 428:38]
  wire [27:0] _GEN_785 = {{27'd0}, _T_3550}; // @[PALU.scala 428:38]
  wire [28:0] _T_3584 = _T_3583 + _GEN_785; // @[PALU.scala 428:38]
  wire [28:0] _GEN_786 = {{28'd0}, _T_3552}; // @[PALU.scala 428:38]
  wire [29:0] _T_3585 = _T_3584 + _GEN_786; // @[PALU.scala 428:38]
  wire [29:0] _GEN_787 = {{29'd0}, _T_3554}; // @[PALU.scala 428:38]
  wire [30:0] _T_3586 = _T_3585 + _GEN_787; // @[PALU.scala 428:38]
  wire [30:0] _GEN_788 = {{30'd0}, _T_3556}; // @[PALU.scala 428:38]
  wire [31:0] _T_3587 = _T_3586 + _GEN_788; // @[PALU.scala 428:38]
  wire [31:0] _T_3589 = _T_3587 - 32'h1; // @[PALU.scala 429:44]
  wire [31:0] _T_3590 = io_in_bits_DecodeIn_data_src2[0] ? _T_3587 : _T_3589; // @[PALU.scala 429:26]
  wire  _T_3593 = io_in_bits_DecodeIn_data_src2[0] ? 1'h0 : io_in_bits_DecodeIn_data_src1[63]; // @[PALU.scala 423:29]
  wire  _T_3595 = io_in_bits_DecodeIn_data_src1[32] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3597 = io_in_bits_DecodeIn_data_src1[33] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3599 = io_in_bits_DecodeIn_data_src1[34] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3601 = io_in_bits_DecodeIn_data_src1[35] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3603 = io_in_bits_DecodeIn_data_src1[36] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3605 = io_in_bits_DecodeIn_data_src1[37] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3607 = io_in_bits_DecodeIn_data_src1[38] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3609 = io_in_bits_DecodeIn_data_src1[39] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3611 = io_in_bits_DecodeIn_data_src1[40] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3613 = io_in_bits_DecodeIn_data_src1[41] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3615 = io_in_bits_DecodeIn_data_src1[42] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3617 = io_in_bits_DecodeIn_data_src1[43] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3619 = io_in_bits_DecodeIn_data_src1[44] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3621 = io_in_bits_DecodeIn_data_src1[45] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3623 = io_in_bits_DecodeIn_data_src1[46] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3625 = io_in_bits_DecodeIn_data_src1[47] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3627 = io_in_bits_DecodeIn_data_src1[48] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3629 = io_in_bits_DecodeIn_data_src1[49] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3631 = io_in_bits_DecodeIn_data_src1[50] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3633 = io_in_bits_DecodeIn_data_src1[51] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3635 = io_in_bits_DecodeIn_data_src1[52] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3637 = io_in_bits_DecodeIn_data_src1[53] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3639 = io_in_bits_DecodeIn_data_src1[54] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3641 = io_in_bits_DecodeIn_data_src1[55] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3643 = io_in_bits_DecodeIn_data_src1[56] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3645 = io_in_bits_DecodeIn_data_src1[57] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3647 = io_in_bits_DecodeIn_data_src1[58] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3649 = io_in_bits_DecodeIn_data_src1[59] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3651 = io_in_bits_DecodeIn_data_src1[60] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3653 = io_in_bits_DecodeIn_data_src1[61] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3655 = io_in_bits_DecodeIn_data_src1[62] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3657 = io_in_bits_DecodeIn_data_src1[63] == _T_3593; // @[PALU.scala 425:59]
  wire  _T_3659 = _T_3655 & _T_3657; // @[PALU.scala 427:113]
  wire  _T_3661 = _T_3653 & (_T_3655 & _T_3657); // @[PALU.scala 427:113]
  wire  _T_3663 = _T_3651 & (_T_3653 & (_T_3655 & _T_3657)); // @[PALU.scala 427:113]
  wire  _T_3665 = _T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))); // @[PALU.scala 427:113]
  wire  _T_3667 = _T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))); // @[PALU.scala 427:113]
  wire  _T_3669 = _T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))); // @[PALU.scala 427:113]
  wire  _T_3671 = _T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))); // @[PALU.scala 427:113]
  wire  _T_3673 = _T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))); // @[PALU.scala 427:113]
  wire  _T_3675 = _T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 &
    _T_3657)))))))); // @[PALU.scala 427:113]
  wire  _T_3677 = _T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (
    _T_3655 & _T_3657))))))))); // @[PALU.scala 427:113]
  wire  _T_3679 = _T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (
    _T_3653 & (_T_3655 & _T_3657)))))))))); // @[PALU.scala 427:113]
  wire  _T_3681 = _T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (
    _T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))); // @[PALU.scala 427:113]
  wire  _T_3683 = _T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (
    _T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))); // @[PALU.scala 427:113]
  wire  _T_3685 = _T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (
    _T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3687 = _T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (
    _T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3689 = _T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (
    _T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3691 = _T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (
    _T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3693 = _T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (
    _T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))
    )))))); // @[PALU.scala 427:113]
  wire  _T_3695 = _T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (
    _T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657
    )))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3697 = _T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (
    _T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (
    _T_3655 & _T_3657))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3699 = _T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (
    _T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (
    _T_3653 & (_T_3655 & _T_3657)))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3701 = _T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (
    _T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (
    _T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3703 = _T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (
    _T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (
    _T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3705 = _T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (
    _T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (
    _T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3707 = _T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (
    _T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (
    _T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3709 = _T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (
    _T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (
    _T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3711 = _T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (_T_3619 & (
    _T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (_T_3639 & (
    _T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657))))))))))))))))))))))
    )))); // @[PALU.scala 427:113]
  wire  _T_3713 = _T_3601 & (_T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (_T_3617 & (
    _T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (_T_3637 & (
    _T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657)))))))))))
    )))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3715 = _T_3599 & (_T_3601 & (_T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (_T_3615 & (
    _T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (_T_3635 & (
    _T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (_T_3655 & _T_3657
    )))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3717 = _T_3597 & (_T_3599 & (_T_3601 & (_T_3603 & (_T_3605 & (_T_3607 & (_T_3609 & (_T_3611 & (_T_3613 & (
    _T_3615 & (_T_3617 & (_T_3619 & (_T_3621 & (_T_3623 & (_T_3625 & (_T_3627 & (_T_3629 & (_T_3631 & (_T_3633 & (
    _T_3635 & (_T_3637 & (_T_3639 & (_T_3641 & (_T_3643 & (_T_3645 & (_T_3647 & (_T_3649 & (_T_3651 & (_T_3653 & (
    _T_3655 & _T_3657))))))))))))))))))))))))))))); // @[PALU.scala 427:113]
  wire  _T_3719 = _T_3595 & _T_3717; // @[PALU.scala 427:113]
  wire [1:0] _T_3720 = _T_3657 + _T_3659; // @[PALU.scala 428:38]
  wire [1:0] _GEN_789 = {{1'd0}, _T_3661}; // @[PALU.scala 428:38]
  wire [2:0] _T_3721 = _T_3720 + _GEN_789; // @[PALU.scala 428:38]
  wire [2:0] _GEN_790 = {{2'd0}, _T_3663}; // @[PALU.scala 428:38]
  wire [3:0] _T_3722 = _T_3721 + _GEN_790; // @[PALU.scala 428:38]
  wire [3:0] _GEN_791 = {{3'd0}, _T_3665}; // @[PALU.scala 428:38]
  wire [4:0] _T_3723 = _T_3722 + _GEN_791; // @[PALU.scala 428:38]
  wire [4:0] _GEN_792 = {{4'd0}, _T_3667}; // @[PALU.scala 428:38]
  wire [5:0] _T_3724 = _T_3723 + _GEN_792; // @[PALU.scala 428:38]
  wire [5:0] _GEN_793 = {{5'd0}, _T_3669}; // @[PALU.scala 428:38]
  wire [6:0] _T_3725 = _T_3724 + _GEN_793; // @[PALU.scala 428:38]
  wire [6:0] _GEN_794 = {{6'd0}, _T_3671}; // @[PALU.scala 428:38]
  wire [7:0] _T_3726 = _T_3725 + _GEN_794; // @[PALU.scala 428:38]
  wire [7:0] _GEN_795 = {{7'd0}, _T_3673}; // @[PALU.scala 428:38]
  wire [8:0] _T_3727 = _T_3726 + _GEN_795; // @[PALU.scala 428:38]
  wire [8:0] _GEN_796 = {{8'd0}, _T_3675}; // @[PALU.scala 428:38]
  wire [9:0] _T_3728 = _T_3727 + _GEN_796; // @[PALU.scala 428:38]
  wire [9:0] _GEN_797 = {{9'd0}, _T_3677}; // @[PALU.scala 428:38]
  wire [10:0] _T_3729 = _T_3728 + _GEN_797; // @[PALU.scala 428:38]
  wire [10:0] _GEN_798 = {{10'd0}, _T_3679}; // @[PALU.scala 428:38]
  wire [11:0] _T_3730 = _T_3729 + _GEN_798; // @[PALU.scala 428:38]
  wire [11:0] _GEN_799 = {{11'd0}, _T_3681}; // @[PALU.scala 428:38]
  wire [12:0] _T_3731 = _T_3730 + _GEN_799; // @[PALU.scala 428:38]
  wire [12:0] _GEN_800 = {{12'd0}, _T_3683}; // @[PALU.scala 428:38]
  wire [13:0] _T_3732 = _T_3731 + _GEN_800; // @[PALU.scala 428:38]
  wire [13:0] _GEN_801 = {{13'd0}, _T_3685}; // @[PALU.scala 428:38]
  wire [14:0] _T_3733 = _T_3732 + _GEN_801; // @[PALU.scala 428:38]
  wire [14:0] _GEN_802 = {{14'd0}, _T_3687}; // @[PALU.scala 428:38]
  wire [15:0] _T_3734 = _T_3733 + _GEN_802; // @[PALU.scala 428:38]
  wire [15:0] _GEN_803 = {{15'd0}, _T_3689}; // @[PALU.scala 428:38]
  wire [16:0] _T_3735 = _T_3734 + _GEN_803; // @[PALU.scala 428:38]
  wire [16:0] _GEN_804 = {{16'd0}, _T_3691}; // @[PALU.scala 428:38]
  wire [17:0] _T_3736 = _T_3735 + _GEN_804; // @[PALU.scala 428:38]
  wire [17:0] _GEN_805 = {{17'd0}, _T_3693}; // @[PALU.scala 428:38]
  wire [18:0] _T_3737 = _T_3736 + _GEN_805; // @[PALU.scala 428:38]
  wire [18:0] _GEN_806 = {{18'd0}, _T_3695}; // @[PALU.scala 428:38]
  wire [19:0] _T_3738 = _T_3737 + _GEN_806; // @[PALU.scala 428:38]
  wire [19:0] _GEN_807 = {{19'd0}, _T_3697}; // @[PALU.scala 428:38]
  wire [20:0] _T_3739 = _T_3738 + _GEN_807; // @[PALU.scala 428:38]
  wire [20:0] _GEN_808 = {{20'd0}, _T_3699}; // @[PALU.scala 428:38]
  wire [21:0] _T_3740 = _T_3739 + _GEN_808; // @[PALU.scala 428:38]
  wire [21:0] _GEN_809 = {{21'd0}, _T_3701}; // @[PALU.scala 428:38]
  wire [22:0] _T_3741 = _T_3740 + _GEN_809; // @[PALU.scala 428:38]
  wire [22:0] _GEN_810 = {{22'd0}, _T_3703}; // @[PALU.scala 428:38]
  wire [23:0] _T_3742 = _T_3741 + _GEN_810; // @[PALU.scala 428:38]
  wire [23:0] _GEN_811 = {{23'd0}, _T_3705}; // @[PALU.scala 428:38]
  wire [24:0] _T_3743 = _T_3742 + _GEN_811; // @[PALU.scala 428:38]
  wire [24:0] _GEN_812 = {{24'd0}, _T_3707}; // @[PALU.scala 428:38]
  wire [25:0] _T_3744 = _T_3743 + _GEN_812; // @[PALU.scala 428:38]
  wire [25:0] _GEN_813 = {{25'd0}, _T_3709}; // @[PALU.scala 428:38]
  wire [26:0] _T_3745 = _T_3744 + _GEN_813; // @[PALU.scala 428:38]
  wire [26:0] _GEN_814 = {{26'd0}, _T_3711}; // @[PALU.scala 428:38]
  wire [27:0] _T_3746 = _T_3745 + _GEN_814; // @[PALU.scala 428:38]
  wire [27:0] _GEN_815 = {{27'd0}, _T_3713}; // @[PALU.scala 428:38]
  wire [28:0] _T_3747 = _T_3746 + _GEN_815; // @[PALU.scala 428:38]
  wire [28:0] _GEN_816 = {{28'd0}, _T_3715}; // @[PALU.scala 428:38]
  wire [29:0] _T_3748 = _T_3747 + _GEN_816; // @[PALU.scala 428:38]
  wire [29:0] _GEN_817 = {{29'd0}, _T_3717}; // @[PALU.scala 428:38]
  wire [30:0] _T_3749 = _T_3748 + _GEN_817; // @[PALU.scala 428:38]
  wire [30:0] _GEN_818 = {{30'd0}, _T_3719}; // @[PALU.scala 428:38]
  wire [31:0] _T_3750 = _T_3749 + _GEN_818; // @[PALU.scala 428:38]
  wire [31:0] _T_3752 = _T_3750 - 32'h1; // @[PALU.scala 429:44]
  wire [31:0] _T_3753 = io_in_bits_DecodeIn_data_src2[0] ? _T_3750 : _T_3752; // @[PALU.scala 429:26]
  wire [63:0] _T_3754 = {_T_3753,_T_3590}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_555 = io_in_bits_Pctrl_isCnt_32 ? _T_3754 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 577:25 579:16]
  wire [63:0] _GEN_556 = io_in_bits_Pctrl_isCnt_8 ? _T_3425 : _GEN_555; // @[PALU.scala 574:24 576:16]
  wire [63:0] cntRes = io_in_bits_Pctrl_isCnt_16 ? _T_3072 : _GEN_556; // @[PALU.scala 571:19 573:16]
  wire [15:0] _GEN_558 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src1[31:16] : 16'h0; // @[PALU.scala 450:37 451:24]
  wire [15:0] _GEN_559 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src2[31:16] : 16'h0; // @[PALU.scala 450:37 452:24]
  wire [15:0] _GEN_560 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src1[31:16] :
    _GEN_558; // @[PALU.scala 447:37 448:24]
  wire [15:0] _GEN_561 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src2[15:0] : _GEN_559
    ; // @[PALU.scala 447:37 449:24]
  wire [15:0] _GEN_562 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src1[15:0] : _GEN_560
    ; // @[PALU.scala 443:37 444:24]
  wire [15:0] _GEN_563 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src2[31:16] :
    _GEN_561; // @[PALU.scala 443:37 445:24]
  wire [15:0] _GEN_564 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src1[15:0] : _GEN_562
    ; // @[PALU.scala 440:31 441:24]
  wire [15:0] _GEN_565 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src2[15:0] : _GEN_563
    ; // @[PALU.scala 440:31 442:24]
  wire [15:0] _GEN_566 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src1[63:48] : 16'h0; // @[PALU.scala 450:37 451:24]
  wire [15:0] _GEN_567 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 ? io_in_bits_DecodeIn_data_src2[63:48] : 16'h0; // @[PALU.scala 450:37 452:24]
  wire [15:0] _GEN_568 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src1[63:48] :
    _GEN_566; // @[PALU.scala 447:37 448:24]
  wire [15:0] _GEN_569 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h3 ? io_in_bits_DecodeIn_data_src2[47:32] :
    _GEN_567; // @[PALU.scala 447:37 449:24]
  wire [15:0] _GEN_570 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src1[47:32] :
    _GEN_568; // @[PALU.scala 443:37 444:24]
  wire [15:0] _GEN_571 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h1 ? io_in_bits_DecodeIn_data_src2[63:48] :
    _GEN_569; // @[PALU.scala 443:37 445:24]
  wire [15:0] _GEN_572 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src1[47:32] :
    _GEN_570; // @[PALU.scala 440:31 441:24]
  wire [15:0] _GEN_573 = io_in_bits_DecodeIn_ctrl_fuOpType[4:3] == 2'h0 ? io_in_bits_DecodeIn_data_src2[47:32] :
    _GEN_571; // @[PALU.scala 440:31 442:24]
  wire [63:0] _T_3841 = {_GEN_572,_GEN_573,_GEN_564,_GEN_565}; // @[Cat.scala 30:58]
  wire [63:0] _T_4012 = {io_in_bits_DecodeIn_data_src1[55:48],io_in_bits_DecodeIn_data_src1[63:56],
    io_in_bits_DecodeIn_data_src1[39:32],io_in_bits_DecodeIn_data_src1[47:40],io_in_bits_DecodeIn_data_src1[23:16],
    io_in_bits_DecodeIn_data_src1[31:24],io_in_bits_DecodeIn_data_src1[7:0],io_in_bits_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_606 = io_in_bits_Pctrl_isSwap_8 ? _T_4012 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 586:25 587:17]
  wire [63:0] swapRes = io_in_bits_Pctrl_isSwap_16 ? _T_3841 : _GEN_606; // @[PALU.scala 584:20 585:17]
  wire [63:0] _GEN_819 = {{32'd0}, io_in_bits_DecodeIn_data_src1[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4016 = _GEN_819 & 64'hffffffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4018 = {io_in_bits_DecodeIn_data_src1[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4020 = _T_4018 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4021 = _T_4016 | _T_4020; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_820 = {{16'd0}, _T_4021[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4026 = _GEN_820 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4028 = {_T_4021[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4030 = _T_4028 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4031 = _T_4026 | _T_4030; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_821 = {{8'd0}, _T_4031[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4036 = _GEN_821 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4038 = {_T_4031[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4040 = _T_4038 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4041 = _T_4036 | _T_4040; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_822 = {{4'd0}, _T_4041[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4046 = _GEN_822 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4048 = {_T_4041[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4050 = _T_4048 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4051 = _T_4046 | _T_4050; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_823 = {{2'd0}, _T_4051[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4056 = _GEN_823 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4058 = {_T_4051[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4060 = _T_4058 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4061 = _T_4056 | _T_4060; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_824 = {{1'd0}, _T_4061[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4066 = _GEN_824 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4068 = {_T_4061[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4070 = _T_4068 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4071 = _T_4066 | _T_4070; // @[Bitwise.scala 103:39]
  wire [63:0] bitrevRes = io_in_bits_Pctrl_isBitrev ? _T_4071 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 592:19 593:19]
  wire  _T_4077 = io_in_bits_DecodeIn_data_src2[0] ? io_in_bits_DecodeIn_data_src1[0] : io_in_bits_DecodeIn_data_src3[0]
    ; // @[PALU.scala 477:46]
  wire  _T_4082 = io_in_bits_DecodeIn_data_src2[1] ? io_in_bits_DecodeIn_data_src1[1] : io_in_bits_DecodeIn_data_src3[1]
    ; // @[PALU.scala 477:46]
  wire  _T_4087 = io_in_bits_DecodeIn_data_src2[2] ? io_in_bits_DecodeIn_data_src1[2] : io_in_bits_DecodeIn_data_src3[2]
    ; // @[PALU.scala 477:46]
  wire  _T_4092 = io_in_bits_DecodeIn_data_src2[3] ? io_in_bits_DecodeIn_data_src1[3] : io_in_bits_DecodeIn_data_src3[3]
    ; // @[PALU.scala 477:46]
  wire  _T_4097 = io_in_bits_DecodeIn_data_src2[4] ? io_in_bits_DecodeIn_data_src1[4] : io_in_bits_DecodeIn_data_src3[4]
    ; // @[PALU.scala 477:46]
  wire  _T_4102 = io_in_bits_DecodeIn_data_src2[5] ? io_in_bits_DecodeIn_data_src1[5] : io_in_bits_DecodeIn_data_src3[5]
    ; // @[PALU.scala 477:46]
  wire  _T_4107 = io_in_bits_DecodeIn_data_src2[6] ? io_in_bits_DecodeIn_data_src1[6] : io_in_bits_DecodeIn_data_src3[6]
    ; // @[PALU.scala 477:46]
  wire  _T_4112 = io_in_bits_DecodeIn_data_src2[7] ? io_in_bits_DecodeIn_data_src1[7] : io_in_bits_DecodeIn_data_src3[7]
    ; // @[PALU.scala 477:46]
  wire  _T_4117 = io_in_bits_DecodeIn_data_src2[8] ? io_in_bits_DecodeIn_data_src1[8] : io_in_bits_DecodeIn_data_src3[8]
    ; // @[PALU.scala 477:46]
  wire  _T_4122 = io_in_bits_DecodeIn_data_src2[9] ? io_in_bits_DecodeIn_data_src1[9] : io_in_bits_DecodeIn_data_src3[9]
    ; // @[PALU.scala 477:46]
  wire  _T_4127 = io_in_bits_DecodeIn_data_src2[10] ? io_in_bits_DecodeIn_data_src1[10] : io_in_bits_DecodeIn_data_src3[
    10]; // @[PALU.scala 477:46]
  wire  _T_4132 = io_in_bits_DecodeIn_data_src2[11] ? io_in_bits_DecodeIn_data_src1[11] : io_in_bits_DecodeIn_data_src3[
    11]; // @[PALU.scala 477:46]
  wire  _T_4137 = io_in_bits_DecodeIn_data_src2[12] ? io_in_bits_DecodeIn_data_src1[12] : io_in_bits_DecodeIn_data_src3[
    12]; // @[PALU.scala 477:46]
  wire  _T_4142 = io_in_bits_DecodeIn_data_src2[13] ? io_in_bits_DecodeIn_data_src1[13] : io_in_bits_DecodeIn_data_src3[
    13]; // @[PALU.scala 477:46]
  wire  _T_4147 = io_in_bits_DecodeIn_data_src2[14] ? io_in_bits_DecodeIn_data_src1[14] : io_in_bits_DecodeIn_data_src3[
    14]; // @[PALU.scala 477:46]
  wire  _T_4152 = io_in_bits_DecodeIn_data_src2[15] ? io_in_bits_DecodeIn_data_src1[15] : io_in_bits_DecodeIn_data_src3[
    15]; // @[PALU.scala 477:46]
  wire  _T_4157 = io_in_bits_DecodeIn_data_src2[16] ? io_in_bits_DecodeIn_data_src1[16] : io_in_bits_DecodeIn_data_src3[
    16]; // @[PALU.scala 477:46]
  wire  _T_4162 = io_in_bits_DecodeIn_data_src2[17] ? io_in_bits_DecodeIn_data_src1[17] : io_in_bits_DecodeIn_data_src3[
    17]; // @[PALU.scala 477:46]
  wire  _T_4167 = io_in_bits_DecodeIn_data_src2[18] ? io_in_bits_DecodeIn_data_src1[18] : io_in_bits_DecodeIn_data_src3[
    18]; // @[PALU.scala 477:46]
  wire  _T_4172 = io_in_bits_DecodeIn_data_src2[19] ? io_in_bits_DecodeIn_data_src1[19] : io_in_bits_DecodeIn_data_src3[
    19]; // @[PALU.scala 477:46]
  wire  _T_4177 = io_in_bits_DecodeIn_data_src2[20] ? io_in_bits_DecodeIn_data_src1[20] : io_in_bits_DecodeIn_data_src3[
    20]; // @[PALU.scala 477:46]
  wire  _T_4182 = io_in_bits_DecodeIn_data_src2[21] ? io_in_bits_DecodeIn_data_src1[21] : io_in_bits_DecodeIn_data_src3[
    21]; // @[PALU.scala 477:46]
  wire  _T_4187 = io_in_bits_DecodeIn_data_src2[22] ? io_in_bits_DecodeIn_data_src1[22] : io_in_bits_DecodeIn_data_src3[
    22]; // @[PALU.scala 477:46]
  wire  _T_4192 = io_in_bits_DecodeIn_data_src2[23] ? io_in_bits_DecodeIn_data_src1[23] : io_in_bits_DecodeIn_data_src3[
    23]; // @[PALU.scala 477:46]
  wire  _T_4197 = io_in_bits_DecodeIn_data_src2[24] ? io_in_bits_DecodeIn_data_src1[24] : io_in_bits_DecodeIn_data_src3[
    24]; // @[PALU.scala 477:46]
  wire  _T_4202 = io_in_bits_DecodeIn_data_src2[25] ? io_in_bits_DecodeIn_data_src1[25] : io_in_bits_DecodeIn_data_src3[
    25]; // @[PALU.scala 477:46]
  wire  _T_4207 = io_in_bits_DecodeIn_data_src2[26] ? io_in_bits_DecodeIn_data_src1[26] : io_in_bits_DecodeIn_data_src3[
    26]; // @[PALU.scala 477:46]
  wire  _T_4212 = io_in_bits_DecodeIn_data_src2[27] ? io_in_bits_DecodeIn_data_src1[27] : io_in_bits_DecodeIn_data_src3[
    27]; // @[PALU.scala 477:46]
  wire  _T_4217 = io_in_bits_DecodeIn_data_src2[28] ? io_in_bits_DecodeIn_data_src1[28] : io_in_bits_DecodeIn_data_src3[
    28]; // @[PALU.scala 477:46]
  wire  _T_4222 = io_in_bits_DecodeIn_data_src2[29] ? io_in_bits_DecodeIn_data_src1[29] : io_in_bits_DecodeIn_data_src3[
    29]; // @[PALU.scala 477:46]
  wire  _T_4227 = io_in_bits_DecodeIn_data_src2[30] ? io_in_bits_DecodeIn_data_src1[30] : io_in_bits_DecodeIn_data_src3[
    30]; // @[PALU.scala 477:46]
  wire  _T_4232 = io_in_bits_DecodeIn_data_src2[31] ? io_in_bits_DecodeIn_data_src1[31] : io_in_bits_DecodeIn_data_src3[
    31]; // @[PALU.scala 477:46]
  wire  _T_4237 = io_in_bits_DecodeIn_data_src2[32] ? io_in_bits_DecodeIn_data_src1[32] : io_in_bits_DecodeIn_data_src3[
    32]; // @[PALU.scala 477:46]
  wire  _T_4242 = io_in_bits_DecodeIn_data_src2[33] ? io_in_bits_DecodeIn_data_src1[33] : io_in_bits_DecodeIn_data_src3[
    33]; // @[PALU.scala 477:46]
  wire  _T_4247 = io_in_bits_DecodeIn_data_src2[34] ? io_in_bits_DecodeIn_data_src1[34] : io_in_bits_DecodeIn_data_src3[
    34]; // @[PALU.scala 477:46]
  wire  _T_4252 = io_in_bits_DecodeIn_data_src2[35] ? io_in_bits_DecodeIn_data_src1[35] : io_in_bits_DecodeIn_data_src3[
    35]; // @[PALU.scala 477:46]
  wire  _T_4257 = io_in_bits_DecodeIn_data_src2[36] ? io_in_bits_DecodeIn_data_src1[36] : io_in_bits_DecodeIn_data_src3[
    36]; // @[PALU.scala 477:46]
  wire  _T_4262 = io_in_bits_DecodeIn_data_src2[37] ? io_in_bits_DecodeIn_data_src1[37] : io_in_bits_DecodeIn_data_src3[
    37]; // @[PALU.scala 477:46]
  wire  _T_4267 = io_in_bits_DecodeIn_data_src2[38] ? io_in_bits_DecodeIn_data_src1[38] : io_in_bits_DecodeIn_data_src3[
    38]; // @[PALU.scala 477:46]
  wire  _T_4272 = io_in_bits_DecodeIn_data_src2[39] ? io_in_bits_DecodeIn_data_src1[39] : io_in_bits_DecodeIn_data_src3[
    39]; // @[PALU.scala 477:46]
  wire  _T_4277 = io_in_bits_DecodeIn_data_src2[40] ? io_in_bits_DecodeIn_data_src1[40] : io_in_bits_DecodeIn_data_src3[
    40]; // @[PALU.scala 477:46]
  wire  _T_4282 = io_in_bits_DecodeIn_data_src2[41] ? io_in_bits_DecodeIn_data_src1[41] : io_in_bits_DecodeIn_data_src3[
    41]; // @[PALU.scala 477:46]
  wire  _T_4287 = io_in_bits_DecodeIn_data_src2[42] ? io_in_bits_DecodeIn_data_src1[42] : io_in_bits_DecodeIn_data_src3[
    42]; // @[PALU.scala 477:46]
  wire  _T_4292 = io_in_bits_DecodeIn_data_src2[43] ? io_in_bits_DecodeIn_data_src1[43] : io_in_bits_DecodeIn_data_src3[
    43]; // @[PALU.scala 477:46]
  wire  _T_4297 = io_in_bits_DecodeIn_data_src2[44] ? io_in_bits_DecodeIn_data_src1[44] : io_in_bits_DecodeIn_data_src3[
    44]; // @[PALU.scala 477:46]
  wire  _T_4302 = io_in_bits_DecodeIn_data_src2[45] ? io_in_bits_DecodeIn_data_src1[45] : io_in_bits_DecodeIn_data_src3[
    45]; // @[PALU.scala 477:46]
  wire  _T_4307 = io_in_bits_DecodeIn_data_src2[46] ? io_in_bits_DecodeIn_data_src1[46] : io_in_bits_DecodeIn_data_src3[
    46]; // @[PALU.scala 477:46]
  wire  _T_4312 = io_in_bits_DecodeIn_data_src2[47] ? io_in_bits_DecodeIn_data_src1[47] : io_in_bits_DecodeIn_data_src3[
    47]; // @[PALU.scala 477:46]
  wire  _T_4317 = io_in_bits_DecodeIn_data_src2[48] ? io_in_bits_DecodeIn_data_src1[48] : io_in_bits_DecodeIn_data_src3[
    48]; // @[PALU.scala 477:46]
  wire  _T_4322 = io_in_bits_DecodeIn_data_src2[49] ? io_in_bits_DecodeIn_data_src1[49] : io_in_bits_DecodeIn_data_src3[
    49]; // @[PALU.scala 477:46]
  wire  _T_4327 = io_in_bits_DecodeIn_data_src2[50] ? io_in_bits_DecodeIn_data_src1[50] : io_in_bits_DecodeIn_data_src3[
    50]; // @[PALU.scala 477:46]
  wire  _T_4332 = io_in_bits_DecodeIn_data_src2[51] ? io_in_bits_DecodeIn_data_src1[51] : io_in_bits_DecodeIn_data_src3[
    51]; // @[PALU.scala 477:46]
  wire  _T_4337 = io_in_bits_DecodeIn_data_src2[52] ? io_in_bits_DecodeIn_data_src1[52] : io_in_bits_DecodeIn_data_src3[
    52]; // @[PALU.scala 477:46]
  wire  _T_4342 = io_in_bits_DecodeIn_data_src2[53] ? io_in_bits_DecodeIn_data_src1[53] : io_in_bits_DecodeIn_data_src3[
    53]; // @[PALU.scala 477:46]
  wire  _T_4347 = io_in_bits_DecodeIn_data_src2[54] ? io_in_bits_DecodeIn_data_src1[54] : io_in_bits_DecodeIn_data_src3[
    54]; // @[PALU.scala 477:46]
  wire  _T_4352 = io_in_bits_DecodeIn_data_src2[55] ? io_in_bits_DecodeIn_data_src1[55] : io_in_bits_DecodeIn_data_src3[
    55]; // @[PALU.scala 477:46]
  wire  _T_4357 = io_in_bits_DecodeIn_data_src2[56] ? io_in_bits_DecodeIn_data_src1[56] : io_in_bits_DecodeIn_data_src3[
    56]; // @[PALU.scala 477:46]
  wire  _T_4362 = io_in_bits_DecodeIn_data_src2[57] ? io_in_bits_DecodeIn_data_src1[57] : io_in_bits_DecodeIn_data_src3[
    57]; // @[PALU.scala 477:46]
  wire  _T_4367 = io_in_bits_DecodeIn_data_src2[58] ? io_in_bits_DecodeIn_data_src1[58] : io_in_bits_DecodeIn_data_src3[
    58]; // @[PALU.scala 477:46]
  wire  _T_4372 = io_in_bits_DecodeIn_data_src2[59] ? io_in_bits_DecodeIn_data_src1[59] : io_in_bits_DecodeIn_data_src3[
    59]; // @[PALU.scala 477:46]
  wire  _T_4377 = io_in_bits_DecodeIn_data_src2[60] ? io_in_bits_DecodeIn_data_src1[60] : io_in_bits_DecodeIn_data_src3[
    60]; // @[PALU.scala 477:46]
  wire  _T_4382 = io_in_bits_DecodeIn_data_src2[61] ? io_in_bits_DecodeIn_data_src1[61] : io_in_bits_DecodeIn_data_src3[
    61]; // @[PALU.scala 477:46]
  wire  _T_4387 = io_in_bits_DecodeIn_data_src2[62] ? io_in_bits_DecodeIn_data_src1[62] : io_in_bits_DecodeIn_data_src3[
    62]; // @[PALU.scala 477:46]
  wire  _T_4392 = io_in_bits_DecodeIn_data_src2[63] ? io_in_bits_DecodeIn_data_src1[63] : io_in_bits_DecodeIn_data_src3[
    63]; // @[PALU.scala 477:46]
  wire [9:0] _T_4401 = {_T_4077,_T_4082,_T_4087,_T_4092,_T_4097,_T_4102,_T_4107,_T_4112,_T_4117,_T_4122}; // @[Cat.scala 30:58]
  wire [18:0] _T_4410 = {_T_4401,_T_4127,_T_4132,_T_4137,_T_4142,_T_4147,_T_4152,_T_4157,_T_4162,_T_4167}; // @[Cat.scala 30:58]
  wire [27:0] _T_4419 = {_T_4410,_T_4172,_T_4177,_T_4182,_T_4187,_T_4192,_T_4197,_T_4202,_T_4207,_T_4212}; // @[Cat.scala 30:58]
  wire [36:0] _T_4428 = {_T_4419,_T_4217,_T_4222,_T_4227,_T_4232,_T_4237,_T_4242,_T_4247,_T_4252,_T_4257}; // @[Cat.scala 30:58]
  wire [45:0] _T_4437 = {_T_4428,_T_4262,_T_4267,_T_4272,_T_4277,_T_4282,_T_4287,_T_4292,_T_4297,_T_4302}; // @[Cat.scala 30:58]
  wire [54:0] _T_4446 = {_T_4437,_T_4307,_T_4312,_T_4317,_T_4322,_T_4327,_T_4332,_T_4337,_T_4342,_T_4347}; // @[Cat.scala 30:58]
  wire [63:0] _T_4455 = {_T_4446,_T_4352,_T_4357,_T_4362,_T_4367,_T_4372,_T_4377,_T_4382,_T_4387,_T_4392}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_825 = {{32'd0}, _T_4455[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4529 = _GEN_825 & 64'hffffffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4531 = {_T_4455[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4533 = _T_4531 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4534 = _T_4529 | _T_4533; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_826 = {{16'd0}, _T_4534[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4539 = _GEN_826 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4541 = {_T_4534[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4543 = _T_4541 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4544 = _T_4539 | _T_4543; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_827 = {{8'd0}, _T_4544[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4549 = _GEN_827 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4551 = {_T_4544[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4553 = _T_4551 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4554 = _T_4549 | _T_4553; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_828 = {{4'd0}, _T_4554[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4559 = _GEN_828 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4561 = {_T_4554[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4563 = _T_4561 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4564 = _T_4559 | _T_4563; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_829 = {{2'd0}, _T_4564[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4569 = _GEN_829 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4571 = {_T_4564[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4573 = _T_4571 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4574 = _T_4569 | _T_4573; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_830 = {{1'd0}, _T_4574[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4579 = _GEN_830 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_4581 = {_T_4574[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_4583 = _T_4581 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] _T_4584 = _T_4579 | _T_4583; // @[Bitwise.scala 103:39]
  wire [63:0] cmixRes = io_in_bits_Pctrl_isCmix ? _T_4584 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 598:17 599:17]
  wire [7:0] _GEN_610 = 3'h0 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[7:0]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_611 = 3'h1 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[15:8]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_612 = 3'h2 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[23:16]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_613 = 3'h3 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[31:24]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_614 = 3'h4 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[39:32]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_615 = 3'h5 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[47:40]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_616 = 3'h6 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[55:48]; // @[PALU.scala 485:31 486:21]
  wire [7:0] _GEN_617 = 3'h7 == io_in_bits_DecodeIn_data_src2[2:0] ? io_in_bits_DecodeIn_data_src1[7:0] :
    io_in_bits_DecodeIn_data_src3[63:56]; // @[PALU.scala 485:31 486:21]
  wire [63:0] _T_4679 = {_GEN_617,_GEN_616,_GEN_615,_GEN_614,_GEN_613,_GEN_612,_GEN_611,_GEN_610}; // @[Cat.scala 30:58]
  wire [63:0] insbRes = io_in_bits_Pctrl_isInsertb ? _T_4679 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 604:20 605:17]
  wire [31:0] _T_4683 = io_in_bits_Pctrl_isPackbb | io_in_bits_Pctrl_isPacktb ? io_in_bits_DecodeIn_data_src2[31:0] :
    io_in_bits_DecodeIn_data_src2[63:32]; // @[PALU.scala 611:25]
  wire [31:0] _T_4687 = io_in_bits_Pctrl_isPackbb | io_in_bits_Pctrl_isPackbt ? io_in_bits_DecodeIn_data_src1[31:0] :
    io_in_bits_DecodeIn_data_src1[63:32]; // @[PALU.scala 612:25]
  wire [63:0] _T_4689 = {_T_4683,_T_4687}; // @[Cat.scala 30:58]
  wire [63:0] _T_4690 = {_T_4687,_T_4683}; // @[Cat.scala 30:58]
  wire [63:0] _T_4691 = io_in_bits_Pctrl_isPackbb | io_in_bits_Pctrl_isPacktt ? _T_4689 : _T_4690; // @[PALU.scala 613:23]
  wire [63:0] packRes = io_in_bits_Pctrl_isPack ? _T_4691 : io_in_bits_DecodeIn_data_src1; // @[PALU.scala 610:17 613:17]
  wire [63:0] _GEN_620 = io_in_bits_Pctrl_isInsertb ? insbRes : adderRes_final; // @[PALU.scala 655:26 656:28 659:28]
  wire  _GEN_621 = io_in_bits_Pctrl_isInsertb ? 1'h0 : adderOV; // @[PALU.scala 655:26 657:39 660:39]
  wire [63:0] _GEN_622 = io_in_bits_Pctrl_isBitrev ? bitrevRes : _GEN_620; // @[PALU.scala 652:25 653:28]
  wire  _GEN_623 = io_in_bits_Pctrl_isBitrev ? 1'h0 : _GEN_621; // @[PALU.scala 652:25 654:39]
  wire [63:0] _GEN_624 = io_in_bits_Pctrl_isPbs ? pbsRes : _GEN_622; // @[PALU.scala 649:22 650:28]
  wire  _GEN_625 = io_in_bits_Pctrl_isPbs ? 1'h0 : _GEN_623; // @[PALU.scala 649:22 651:39]
  wire [63:0] _GEN_626 = io_in_bits_Pctrl_isUnpack ? unpackRes : _GEN_624; // @[PALU.scala 646:25 647:28]
  wire  _GEN_627 = io_in_bits_Pctrl_isUnpack ? 1'h0 : _GEN_625; // @[PALU.scala 646:25 648:39]
  wire [63:0] _GEN_628 = io_in_bits_Pctrl_isCnt ? cntRes : _GEN_626; // @[PALU.scala 643:22 644:28]
  wire  _GEN_629 = io_in_bits_Pctrl_isCnt ? 1'h0 : _GEN_627; // @[PALU.scala 643:22 645:39]
  wire [63:0] _GEN_630 = io_in_bits_Pctrl_isSat ? satRes : _GEN_628; // @[PALU.scala 640:22 641:28]
  wire  _GEN_631 = io_in_bits_Pctrl_isSat ? satOV : _GEN_629; // @[PALU.scala 640:22 642:39]
  wire [63:0] _GEN_632 = io_in_bits_Pctrl_isClip ? clipRes : _GEN_630; // @[PALU.scala 637:23 638:28]
  wire  _GEN_633 = io_in_bits_Pctrl_isClip ? clipOV : _GEN_631; // @[PALU.scala 637:23 639:39]
  wire [63:0] _GEN_634 = io_in_bits_Pctrl_isCompare ? compareRes : _GEN_632; // @[PALU.scala 634:26 635:28]
  wire  _GEN_635 = io_in_bits_Pctrl_isCompare ? 1'h0 : _GEN_633; // @[PALU.scala 634:26 636:39]
  wire [63:0] _GEN_636 = io_in_bits_Pctrl_isShifter ? shifterRes : _GEN_634; // @[PALU.scala 631:26 632:28]
  wire  _GEN_637 = io_in_bits_Pctrl_isShifter ? shifterOV : _GEN_635; // @[PALU.scala 631:26 633:39]
  wire [63:0] _GEN_638 = io_in_bits_Pctrl_isAdder ? adderRes_final : _GEN_636; // @[PALU.scala 628:24 629:28]
  wire  _GEN_639 = io_in_bits_Pctrl_isAdder ? adderOV : _GEN_637; // @[PALU.scala 628:24 630:39]
  wire [63:0] _GEN_640 = io_in_bits_Pctrl_isCmix ? cmixRes : _GEN_638; // @[PALU.scala 625:23 626:28]
  wire  _GEN_641 = io_in_bits_Pctrl_isCmix ? 1'h0 : _GEN_639; // @[PALU.scala 625:23 627:39]
  wire [63:0] _GEN_642 = io_in_bits_Pctrl_isSwap ? swapRes : _GEN_640; // @[PALU.scala 622:23 623:28]
  wire  _GEN_643 = io_in_bits_Pctrl_isSwap ? 1'h0 : _GEN_641; // @[PALU.scala 622:23 624:39]
  wire [63:0] _GEN_644 = io_in_bits_Pctrl_isMaxMin ? maxminRes : _GEN_642; // @[PALU.scala 619:25 620:28]
  wire  _GEN_645 = io_in_bits_Pctrl_isMaxMin ? 1'h0 : _GEN_643; // @[PALU.scala 619:25 621:39]
  assign io_in_ready = ~io_in_valid | _T_1; // @[PALU.scala 37:27]
  assign io_out_valid = io_in_valid; // @[PALU.scala 38:17]
  assign io_out_bits_result = io_in_bits_Pctrl_isPack ? packRes : _GEN_644; // @[PALU.scala 616:17 617:28]
  assign io_out_bits_DecodeOut_cf_pc = io_in_bits_DecodeIn_cf_pc; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_cf_runahead_checkpoint_id = io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_ctrl_rfWen = io_in_bits_DecodeIn_ctrl_rfWen; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_ctrl_rfDest = io_in_bits_DecodeIn_ctrl_rfDest; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_pext_OV = io_in_bits_Pctrl_isPack ? 1'h0 : _GEN_645; // @[PALU.scala 616:17 618:39]
  assign io_out_bits_DecodeOut_InstNo = io_in_bits_DecodeIn_InstNo; // @[PALU.scala 39:27]
  assign io_out_bits_DecodeOut_InstFlag = io_in_bits_DecodeIn_InstFlag; // @[PALU.scala 39:27]
endmodule
module PMDU_1(
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_DecodeIn_cf_pc,
  input  [63:0]  io_in_bits_DecodeIn_cf_runahead_checkpoint_id,
  input  [6:0]   io_in_bits_DecodeIn_ctrl_fuOpType,
  input          io_in_bits_DecodeIn_ctrl_rfWen,
  input  [4:0]   io_in_bits_DecodeIn_ctrl_rfDest,
  input  [63:0]  io_in_bits_DecodeIn_data_src1,
  input  [63:0]  io_in_bits_DecodeIn_data_src2,
  input  [63:0]  io_in_bits_DecodeIn_data_src3,
  input  [4:0]   io_in_bits_DecodeIn_InstNo,
  input          io_in_bits_DecodeIn_InstFlag,
  input          io_in_bits_Pctrl_isMul_16,
  input          io_in_bits_Pctrl_isMul_8,
  input          io_in_bits_Pctrl_isMSW_3232,
  input          io_in_bits_Pctrl_isMSW_3216,
  input          io_in_bits_Pctrl_isS1632,
  input          io_in_bits_Pctrl_isS1664,
  input          io_in_bits_Pctrl_is832,
  input          io_in_bits_Pctrl_is3264,
  input          io_in_bits_Pctrl_is1664,
  input          io_in_bits_Pctrl_isQ15orQ31,
  input          io_in_bits_Pctrl_isC31,
  input          io_in_bits_Pctrl_isQ15_64ONLY,
  input          io_in_bits_Pctrl_isQ63_64ONLY,
  input          io_in_bits_Pctrl_isMul_32_64ONLY,
  input          io_in_bits_Pctrl_isPMA_64ONLY,
  input  [17:0]  io_in_bits_Pctrl_mulres9_0,
  input  [17:0]  io_in_bits_Pctrl_mulres9_1,
  input  [17:0]  io_in_bits_Pctrl_mulres9_2,
  input  [17:0]  io_in_bits_Pctrl_mulres9_3,
  input  [33:0]  io_in_bits_Pctrl_mulres17_0,
  input  [33:0]  io_in_bits_Pctrl_mulres17_1,
  input  [65:0]  io_in_bits_Pctrl_mulres33_0,
  input  [129:0] io_in_bits_Pctrl_mulres65_0,
  input          io_out_ready,
  output         io_out_valid,
  output [63:0]  io_out_bits_result,
  output [38:0]  io_out_bits_DecodeOut_cf_pc,
  output [63:0]  io_out_bits_DecodeOut_cf_runahead_checkpoint_id,
  output [6:0]   io_out_bits_DecodeOut_ctrl_fuOpType,
  output         io_out_bits_DecodeOut_ctrl_rfWen,
  output [4:0]   io_out_bits_DecodeOut_ctrl_rfDest,
  output [63:0]  io_out_bits_DecodeOut_data_src1,
  output [63:0]  io_out_bits_DecodeOut_data_src2,
  output [63:0]  io_out_bits_DecodeOut_data_src3,
  output         io_out_bits_DecodeOut_pext_OV,
  output [4:0]   io_out_bits_DecodeOut_InstNo,
  output         io_out_bits_DecodeOut_InstFlag,
  output         io_FirstStageFire
);
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [32:0] _T_718 = {io_out_bits_DecodeOut_data_src3[63],io_out_bits_DecodeOut_data_src3[63:32]}; // @[Cat.scala 30:58]
  wire [1:0] _T_1035 = io_out_bits_DecodeOut_data_src3[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1036 = {_T_1035,io_out_bits_DecodeOut_data_src3[63:32]}; // @[Cat.scala 30:58]
  wire  _T_467 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h4; // @[PMDU.scala 849:59]
  wire [31:0] _T_469 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h4 ? io_out_bits_DecodeOut_data_src3[63:32] : 32'h0
    ; // @[PMDU.scala 849:45]
  wire [32:0] _T_471 = {_T_469[31],_T_469}; // @[Cat.scala 30:58]
  wire [33:0] _GEN_88 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _T_471} : 34'h0; // @[PMDU.scala 836:50 865:34]
  wire [33:0] _GEN_101 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_88; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_113 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_101; // @[PMDU.scala 735:40]
  wire [33:0] _GEN_223 = io_in_bits_Pctrl_is832 ? {{2'd0}, io_out_bits_DecodeOut_data_src3[63:32]} : _GEN_113; // @[PMDU.scala 1051:39 1078:30]
  wire [33:0] _GEN_244 = io_in_bits_Pctrl_isS1664 ? _GEN_113 : _GEN_223; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_257 = io_in_bits_Pctrl_isS1632 ? _T_1036 : _GEN_244; // @[PMDU.scala 1000:41 1020:30]
  wire [33:0] _GEN_273 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_718} : _GEN_257; // @[PMDU.scala 963:44 979:30]
  wire [33:0] adder34_0_1 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_718} : _GEN_273; // @[PMDU.scala 929:38 938:30]
  wire [32:0] _T_638 = {io_out_bits_DecodeOut_data_src3[31],io_out_bits_DecodeOut_data_src3[31:0]}; // @[Cat.scala 30:58]
  wire [1:0] _T_968 = io_out_bits_DecodeOut_data_src3[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_969 = {_T_968,io_out_bits_DecodeOut_data_src3[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_417 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h4 ? io_out_bits_DecodeOut_data_src3[31:0] : 32'h0; // @[PMDU.scala 849:45]
  wire [32:0] _T_419 = {_T_417[31],_T_417}; // @[Cat.scala 30:58]
  wire [33:0] _GEN_85 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _T_419} : 34'h0; // @[PMDU.scala 836:50 865:34]
  wire [33:0] _GEN_98 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_85; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_110 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_98; // @[PMDU.scala 735:40]
  wire [33:0] _GEN_218 = io_in_bits_Pctrl_is832 ? {{2'd0}, io_out_bits_DecodeOut_data_src3[31:0]} : _GEN_110; // @[PMDU.scala 1051:39 1078:30]
  wire [33:0] _GEN_239 = io_in_bits_Pctrl_isS1664 ? _GEN_110 : _GEN_218; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_252 = io_in_bits_Pctrl_isS1632 ? _T_969 : _GEN_239; // @[PMDU.scala 1000:41 1020:30]
  wire [33:0] _GEN_270 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_638} : _GEN_252; // @[PMDU.scala 963:44 979:30]
  wire [33:0] adder34_0_0 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_638} : _GEN_270; // @[PMDU.scala 929:38 938:30]
  wire [70:0] _T_12 = {adder34_0_1,3'h0,adder34_0_0}; // @[Cat.scala 30:58]
  wire [64:0] _T_512 = {io_out_bits_DecodeOut_data_src3[63],io_out_bits_DecodeOut_data_src3}; // @[Cat.scala 30:58]
  wire  _T_533 = ~(_T_467 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h1d); // @[PMDU.scala 904:31]
  wire [1:0] _T_555 = io_out_bits_DecodeOut_data_src3[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_556 = {_T_555,io_out_bits_DecodeOut_data_src3}; // @[Cat.scala 30:58]
  wire [65:0] _T_557 = _T_533 ? _T_556 : 66'h0; // @[PMDU.scala 908:33]
  wire [70:0] _GEN_66 = io_in_bits_Pctrl_isPMA_64ONLY ? {{5'd0}, _T_557} : _T_12; // @[PMDU.scala 728:15 902:50 908:27]
  wire [70:0] _GEN_72 = io_in_bits_Pctrl_isQ63_64ONLY ? {{6'd0}, _T_512} : _GEN_66; // @[PMDU.scala 886:50 888:27]
  wire [70:0] _GEN_79 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_12 : _GEN_72; // @[PMDU.scala 728:15 884:53]
  wire [70:0] _GEN_92 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_12 : _GEN_79; // @[PMDU.scala 728:15 836:50]
  wire [70:0] _GEN_104 = io_in_bits_Pctrl_isMul_8 ? _T_12 : _GEN_92; // @[PMDU.scala 728:15 779:45]
  wire [70:0] _GEN_116 = io_in_bits_Pctrl_isMul_16 ? _T_12 : _GEN_104; // @[PMDU.scala 728:15 735:40]
  wire  _T_1198 = ~io_out_bits_DecodeOut_ctrl_fuOpType[4]; // @[PMDU.scala 1090:24]
  wire [65:0] _T_1216 = {2'h0,io_out_bits_DecodeOut_data_src3}; // @[Cat.scala 30:58]
  wire [65:0] _GEN_176 = _T_1198 ? _T_556 : _T_1216; // @[PMDU.scala 676:24 677:15 679:15]
  wire [31:0] _T_1413 = io_out_bits_DecodeOut_ctrl_fuOpType[4] ? 32'h0 : io_out_bits_DecodeOut_data_src3[31:0]; // @[PMDU.scala 1186:29]
  wire [70:0] _GEN_195 = io_in_bits_Pctrl_isC31 ? {{39'd0}, _T_1413} : _GEN_116; // @[PMDU.scala 1183:39 1186:23]
  wire [70:0] _GEN_200 = io_in_bits_Pctrl_isQ15orQ31 ? {{38'd0}, _T_638} : _GEN_195; // @[PMDU.scala 1149:44 1167:23]
  wire [70:0] _GEN_204 = io_in_bits_Pctrl_is1664 ? {{7'd0}, io_out_bits_DecodeOut_data_src3} : _GEN_200; // @[PMDU.scala 1126:40 1136:23]
  wire [70:0] _GEN_211 = io_in_bits_Pctrl_is3264 ? {{5'd0}, _GEN_176} : _GEN_204; // @[PMDU.scala 1089:40 1098:23]
  wire [70:0] _GEN_229 = io_in_bits_Pctrl_is832 ? _GEN_116 : _GEN_211; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_235 = io_in_bits_Pctrl_isS1664 ? {{7'd0}, io_out_bits_DecodeOut_data_src1} : _GEN_229; // @[PMDU.scala 1046:41 1047:19]
  wire [70:0] _GEN_262 = io_in_bits_Pctrl_isS1632 ? _GEN_116 : _GEN_235; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_279 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_116 : _GEN_262; // @[PMDU.scala 963:44]
  wire [70:0] adder68_0 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_116 : _GEN_279; // @[PMDU.scala 929:38]
  wire  _T_686 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h1; // @[PMDU.scala 933:69]
  wire  _T_687 = io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h2 & io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h1; // @[PMDU.scala 933:52]
  wire [32:0] _T_720 = _T_687 ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire  _T_694 = io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h3; // @[PMDU.scala 935:40]
  wire  _T_697 = io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h3 & _T_686; // @[PMDU.scala 935:52]
  wire [32:0] _T_703 = io_in_bits_Pctrl_mulres65_0[63:31] + 33'h1; // @[PMDU.scala 936:164]
  wire [32:0] _T_705 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_703 : io_in_bits_Pctrl_mulres65_0[63:31]; // @[PMDU.scala 936:41]
  wire [33:0] _T_711 = io_in_bits_Pctrl_mulres65_0[63:30] + 34'h1; // @[PMDU.scala 937:164]
  wire [33:0] _T_713 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_711 : io_in_bits_Pctrl_mulres65_0[63:30]; // @[PMDU.scala 937:41]
  wire [31:0] _T_715 = ~_T_697 ? _T_705[32:1] : _T_713[32:1]; // @[PMDU.scala 936:32]
  wire [32:0] _T_722 = {_T_715[31],_T_715}; // @[Cat.scala 30:58]
  wire [32:0] _T_723 = _T_720 ^ _T_722; // @[PMDU.scala 939:53]
  wire  _T_847 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h7; // @[PMDU.scala 968:41]
  wire  _T_880 = io_out_bits_DecodeOut_data_src1[63:32] == 32'h80000000; // @[PMDU.scala 975:62]
  wire  _T_855 = _T_694 | io_out_bits_DecodeOut_ctrl_fuOpType[6:4] == 3'h5 | io_out_bits_DecodeOut_ctrl_fuOpType[6:4]
     == 3'h7; // @[PMDU.scala 969:93]
  wire [15:0] _T_858 = _T_855 ? io_out_bits_DecodeOut_data_src2[63:48] : io_out_bits_DecodeOut_data_src2[47:32]; // @[PMDU.scala 970:36]
  wire [32:0] _T_864 = io_in_bits_Pctrl_mulres65_0[47:15] + 33'h1; // @[PMDU.scala 971:165]
  wire [32:0] _T_866 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_864 : io_in_bits_Pctrl_mulres65_0[47:15]; // @[PMDU.scala 971:42]
  wire [32:0] _T_872 = io_in_bits_Pctrl_mulres65_0[46:14] + 33'h1; // @[PMDU.scala 972:164]
  wire [32:0] _T_874 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_872 : io_in_bits_Pctrl_mulres65_0[46:14]; // @[PMDU.scala 972:41]
  wire [31:0] _T_876 = ~_T_847 ? _T_866[32:1] : _T_874[32:1]; // @[PMDU.scala 971:33]
  wire [31:0] _GEN_146 = _T_847 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80000000 & _T_858 == 16'h8000 ? 32'h7fffffff
     : _T_876; // @[PMDU.scala 975:127 974:23 977:27]
  wire [32:0] _T_892 = {_GEN_146[31],_GEN_146}; // @[Cat.scala 30:58]
  wire  _T_934 = io_out_bits_DecodeOut_ctrl_fuOpType[6:1] == 6'h13; // @[PMDU.scala 1002:95]
  wire  _T_935 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h34 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h36 |
    io_out_bits_DecodeOut_ctrl_fuOpType[6:1] == 6'h13; // @[PMDU.scala 1002:78]
  wire [33:0] _T_1038 = _T_935 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_1041 = io_in_bits_Pctrl_mulres65_0[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1042 = {_T_1041,io_in_bits_Pctrl_mulres65_0[31:0]}; // @[Cat.scala 30:58]
  wire [33:0] _T_1043 = _T_1038 ^ _T_1042; // @[PMDU.scala 1021:57]
  wire  _T_402 = io_out_bits_DecodeOut_ctrl_fuOpType[4:3] == 2'h1; // @[PMDU.scala 838:40]
  wire  _T_404 = io_out_bits_DecodeOut_ctrl_fuOpType[4:3] == 2'h2; // @[PMDU.scala 839:40]
  wire [15:0] _T_460 = _T_404 ? io_out_bits_DecodeOut_data_src1[47:32] : io_out_bits_DecodeOut_data_src1[63:48]; // @[PMDU.scala 842:70]
  wire [15:0] _T_461 = _T_402 ? io_out_bits_DecodeOut_data_src1[47:32] : _T_460; // @[PMDU.scala 842:40]
  wire [15:0] _T_464 = _T_402 ? io_out_bits_DecodeOut_data_src2[47:32] : io_out_bits_DecodeOut_data_src2[63:48]; // @[PMDU.scala 843:40]
  wire  _T_476 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h6; // @[PMDU.scala 853:44]
  wire [30:0] _GEN_49 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h6 ? 31'h7fff : 31'h7fffffff; // @[PMDU.scala 853:57 854:36 856:36]
  wire [16:0] _T_482 = io_in_bits_Pctrl_mulres65_0[30] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_483 = {_T_482,io_in_bits_Pctrl_mulres65_0[30:15]}; // @[Cat.scala 30:58]
  wire [32:0] _T_485 = {io_in_bits_Pctrl_mulres65_0[31],io_in_bits_Pctrl_mulres65_0[31:0]}; // @[Cat.scala 30:58]
  wire [33:0] _T_486 = {_T_485, 1'h0}; // @[PMDU.scala 862:64]
  wire [32:0] _T_489 = {_T_486[31],_T_486[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_50 = _T_476 ? _T_483 : _T_489; // @[PMDU.scala 859:57 860:36 862:36]
  wire [32:0] _GEN_52 = _T_461 == 16'h8000 & _T_464 == 16'h8000 ? {{2'd0}, _GEN_49} : _GEN_50; // @[PMDU.scala 851:77]
  wire [33:0] _GEN_89 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _GEN_52} : 34'h0; // @[PMDU.scala 836:50 866:34]
  wire [33:0] _GEN_102 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_89; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_114 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_102; // @[PMDU.scala 735:40]
  wire  _T_1156 = ~_T_476; // @[PMDU.scala 1073:38]
  wire [14:0] _T_1160 = io_in_bits_Pctrl_mulres17_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1161 = {_T_1160,io_in_bits_Pctrl_mulres17_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1162 = {15'h0,io_in_bits_Pctrl_mulres17_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_170 = _T_1156 ? _T_1161 : _T_1162; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_224 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_170} : _GEN_114; // @[PMDU.scala 1051:39 1079:30]
  wire [33:0] _GEN_245 = io_in_bits_Pctrl_isS1664 ? _GEN_114 : _GEN_224; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_258 = io_in_bits_Pctrl_isS1632 ? _T_1043 : _GEN_245; // @[PMDU.scala 1000:41 1021:30]
  wire [33:0] _GEN_274 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_892} : _GEN_258; // @[PMDU.scala 963:44 980:30]
  wire [33:0] adder34_1_1 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_723} : _GEN_274; // @[PMDU.scala 929:38 939:30]
  wire [32:0] _T_623 = io_in_bits_Pctrl_mulres33_0[63:31] + 33'h1; // @[PMDU.scala 936:120]
  wire [32:0] _T_625 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_623 : io_in_bits_Pctrl_mulres33_0[63:31]; // @[PMDU.scala 936:41]
  wire [33:0] _T_631 = io_in_bits_Pctrl_mulres33_0[63:30] + 34'h1; // @[PMDU.scala 937:120]
  wire [33:0] _T_633 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_631 : io_in_bits_Pctrl_mulres33_0[63:30]; // @[PMDU.scala 937:41]
  wire [31:0] _T_635 = ~_T_697 ? _T_625[32:1] : _T_633[32:1]; // @[PMDU.scala 936:32]
  wire [32:0] _T_642 = {_T_635[31],_T_635}; // @[Cat.scala 30:58]
  wire [32:0] _T_643 = _T_720 ^ _T_642; // @[PMDU.scala 939:53]
  wire  _T_803 = io_out_bits_DecodeOut_data_src1[31:0] == 32'h80000000; // @[PMDU.scala 975:62]
  wire [15:0] _T_781 = _T_855 ? io_out_bits_DecodeOut_data_src2[31:16] : io_out_bits_DecodeOut_data_src2[15:0]; // @[PMDU.scala 970:36]
  wire [32:0] _T_787 = io_in_bits_Pctrl_mulres33_0[47:15] + 33'h1; // @[PMDU.scala 971:121]
  wire [32:0] _T_789 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_787 : io_in_bits_Pctrl_mulres33_0[47:15]; // @[PMDU.scala 971:42]
  wire [32:0] _T_795 = io_in_bits_Pctrl_mulres33_0[46:14] + 33'h1; // @[PMDU.scala 972:120]
  wire [32:0] _T_797 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _T_795 : io_in_bits_Pctrl_mulres33_0[46:14]; // @[PMDU.scala 972:41]
  wire [31:0] _T_799 = ~_T_847 ? _T_789[32:1] : _T_797[32:1]; // @[PMDU.scala 971:33]
  wire [31:0] _GEN_139 = _T_847 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80000000 & _T_781 == 16'h8000 ? 32'h7fffffff
     : _T_799; // @[PMDU.scala 975:127 974:23 977:27]
  wire [32:0] _T_815 = {_GEN_139[31],_GEN_139}; // @[Cat.scala 30:58]
  wire  _T_922 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h5; // @[PMDU.scala 1001:61]
  wire  _T_924 = io_out_bits_DecodeOut_ctrl_fuOpType[6:5] == 2'h1; // @[PMDU.scala 1001:91]
  wire  _T_929 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] < 4'h3 | io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h5 &
    io_out_bits_DecodeOut_ctrl_fuOpType[6:5] == 2'h1 & io_out_bits_DecodeOut_ctrl_fuOpType[4:3] != 2'h0; // @[PMDU.scala 1001:44]
  wire [31:0] _T_962 = _T_929 ? io_in_bits_Pctrl_mulres33_0[31:0] : io_in_bits_Pctrl_mulres17_1[31:0]; // @[PMDU.scala 1011:39]
  wire [1:0] _T_974 = _T_962[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_975 = {_T_974,_T_962}; // @[Cat.scala 30:58]
  wire [33:0] _T_976 = _T_1038 ^ _T_975; // @[PMDU.scala 1021:57]
  wire [15:0] _T_408 = _T_404 ? io_out_bits_DecodeOut_data_src1[15:0] : io_out_bits_DecodeOut_data_src1[31:16]; // @[PMDU.scala 842:70]
  wire [15:0] _T_409 = _T_402 ? io_out_bits_DecodeOut_data_src1[15:0] : _T_408; // @[PMDU.scala 842:40]
  wire [15:0] _T_412 = _T_402 ? io_out_bits_DecodeOut_data_src2[15:0] : io_out_bits_DecodeOut_data_src2[31:16]; // @[PMDU.scala 843:40]
  wire  _T_422 = _T_409 == 16'h8000 & _T_412 == 16'h8000; // @[PMDU.scala 851:50]
  wire [16:0] _T_430 = io_in_bits_Pctrl_mulres33_0[30] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_431 = {_T_430,io_in_bits_Pctrl_mulres33_0[30:15]}; // @[Cat.scala 30:58]
  wire [32:0] _T_433 = {io_in_bits_Pctrl_mulres33_0[31],io_in_bits_Pctrl_mulres33_0[31:0]}; // @[Cat.scala 30:58]
  wire [33:0] _T_434 = {_T_433, 1'h0}; // @[PMDU.scala 862:64]
  wire [32:0] _T_437 = {_T_434[31],_T_434[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_41 = _T_476 ? _T_431 : _T_437; // @[PMDU.scala 859:57 860:36 862:36]
  wire [32:0] _GEN_43 = _T_409 == 16'h8000 & _T_412 == 16'h8000 ? {{2'd0}, _GEN_49} : _GEN_41; // @[PMDU.scala 851:77]
  wire [33:0] _GEN_86 = io_in_bits_Pctrl_isQ15_64ONLY ? {{1'd0}, _GEN_43} : 34'h0; // @[PMDU.scala 836:50 866:34]
  wire [33:0] _GEN_99 = io_in_bits_Pctrl_isMul_8 ? 34'h0 : _GEN_86; // @[PMDU.scala 779:45]
  wire [33:0] _GEN_111 = io_in_bits_Pctrl_isMul_16 ? 34'h0 : _GEN_99; // @[PMDU.scala 735:40]
  wire [14:0] _T_1121 = io_in_bits_Pctrl_mulres9_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1122 = {_T_1121,io_in_bits_Pctrl_mulres9_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1123 = {15'h0,io_in_bits_Pctrl_mulres9_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_166 = _T_1156 ? _T_1122 : _T_1123; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_219 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_166} : _GEN_111; // @[PMDU.scala 1051:39 1079:30]
  wire [33:0] _GEN_240 = io_in_bits_Pctrl_isS1664 ? _GEN_111 : _GEN_219; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_253 = io_in_bits_Pctrl_isS1632 ? _T_976 : _GEN_240; // @[PMDU.scala 1000:41 1021:30]
  wire [33:0] _GEN_271 = io_in_bits_Pctrl_isMSW_3216 ? {{1'd0}, _T_815} : _GEN_253; // @[PMDU.scala 963:44 980:30]
  wire [33:0] adder34_1_0 = io_in_bits_Pctrl_isMSW_3232 ? {{1'd0}, _T_643} : _GEN_271; // @[PMDU.scala 929:38 939:30]
  wire [70:0] _T_13 = {adder34_1_1,3'h0,adder34_1_0}; // @[Cat.scala 30:58]
  wire [64:0] _T_515 = {io_in_bits_Pctrl_mulres65_0[63],io_in_bits_Pctrl_mulres65_0[63:0]}; // @[Cat.scala 30:58]
  wire  _T_538 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h5 | io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h7; // @[PMDU.scala 905:59]
  wire  _T_541 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h5 | io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h7 |
    _T_934; // @[PMDU.scala 905:90]
  wire [65:0] _T_559 = _T_541 ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_563 = io_in_bits_Pctrl_mulres33_0[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_564 = {_T_563,io_in_bits_Pctrl_mulres33_0[63:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_565 = _T_559 ^ _T_564; // @[PMDU.scala 909:47]
  wire [70:0] _GEN_67 = io_in_bits_Pctrl_isPMA_64ONLY ? {{5'd0}, _T_565} : _T_13; // @[PMDU.scala 729:15 902:50 909:27]
  wire [70:0] _GEN_73 = io_in_bits_Pctrl_isQ63_64ONLY ? {{6'd0}, _T_515} : _GEN_67; // @[PMDU.scala 886:50 889:27]
  wire [70:0] _GEN_80 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_13 : _GEN_73; // @[PMDU.scala 729:15 884:53]
  wire [70:0] _GEN_93 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_13 : _GEN_80; // @[PMDU.scala 729:15 836:50]
  wire [70:0] _GEN_105 = io_in_bits_Pctrl_isMul_8 ? _T_13 : _GEN_93; // @[PMDU.scala 729:15 779:45]
  wire [70:0] _GEN_117 = io_in_bits_Pctrl_isMul_16 ? _T_13 : _GEN_105; // @[PMDU.scala 729:15 735:40]
  wire [31:0] _T_1107 = io_in_bits_Pctrl_mulres65_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1108 = {_T_1107,io_in_bits_Pctrl_mulres65_0[31:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1218 = io_out_bits_DecodeOut_ctrl_fuOpType[0] ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_1205 = {io_in_bits_Pctrl_mulres33_0[64],io_in_bits_Pctrl_mulres33_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1206 = {1'h0,io_in_bits_Pctrl_mulres33_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _GEN_174 = _T_1198 ? _T_1205 : _T_1206; // @[PMDU.scala 676:24 677:15 679:15]
  wire [65:0] _T_1219 = _T_1218 ^ _GEN_174; // @[PMDU.scala 1099:41]
  wire  _T_1258 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h56; // @[PMDU.scala 1128:90]
  wire  _T_1260 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h5e; // @[PMDU.scala 1128:119]
  wire  _T_1261 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h45 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h55 |
    io_out_bits_DecodeOut_ctrl_fuOpType == 7'h56 | io_out_bits_DecodeOut_ctrl_fuOpType == 7'h5e; // @[PMDU.scala 1128:107]
  wire [63:0] _T_1279 = _T_1261 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1269 = _T_467 ? io_in_bits_Pctrl_mulres33_0[31:0] : io_in_bits_Pctrl_mulres17_0[31:0]; // @[PMDU.scala 1132:23]
  wire [31:0] _T_1282 = _T_1269[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1283 = {_T_1282,_T_1269}; // @[Cat.scala 30:58]
  wire [63:0] _T_1284 = _T_1279 ^ _T_1283; // @[PMDU.scala 1137:50]
  wire [1:0] _T_1285 = {_T_1261,1'h0}; // @[Cat.scala 30:58]
  wire  _T_1266 = io_out_bits_DecodeOut_ctrl_fuOpType == 7'h4d | _T_1258 | _T_1260; // @[PMDU.scala 1129:78]
  wire [1:0] _T_1286 = {_T_1266,1'h0}; // @[Cat.scala 30:58]
  wire [2:0] _T_1287 = _T_1285 + _T_1286; // @[PMDU.scala 1137:101]
  wire [63:0] _GEN_303 = {{61'd0}, _T_1287}; // @[PMDU.scala 1137:69]
  wire [63:0] _T_1289 = _T_1284 + _GEN_303; // @[PMDU.scala 1137:69]
  wire  _T_1344 = _T_686 ? _T_402 : io_out_bits_DecodeOut_ctrl_fuOpType[4:3] == 2'h0; // @[PMDU.scala 1154:25]
  wire  _T_1349 = _T_686 ? _T_404 : _T_402; // @[PMDU.scala 1155:25]
  wire [15:0] _T_1353 = _T_1349 ? io_out_bits_DecodeOut_data_src1[15:0] : io_out_bits_DecodeOut_data_src1[31:16]; // @[PMDU.scala 1156:55]
  wire [15:0] _T_1354 = _T_1344 ? io_out_bits_DecodeOut_data_src1[15:0] : _T_1353; // @[PMDU.scala 1156:33]
  wire [15:0] _T_1357 = _T_1344 ? io_out_bits_DecodeOut_data_src2[15:0] : io_out_bits_DecodeOut_data_src2[31:16]; // @[PMDU.scala 1157:33]
  wire [63:0] _T_1364 = _T_476 ? 64'h7fff : 64'h7fffffff; // @[PMDU.scala 1163:28]
  wire [31:0] _T_1365 = io_in_bits_Pctrl_mulres65_0[31:0]; // @[PMDU.scala 1165:48]
  wire [16:0] _T_1367 = _T_1365[31:15]; // @[PMDU.scala 1165:62]
  wire [46:0] _T_1370 = _T_1367[16] ? 47'h7fffffffffff : 47'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1371 = {_T_1370,_T_1367}; // @[Cat.scala 30:58]
  wire [32:0] _T_1372 = {io_in_bits_Pctrl_mulres65_0[31:0], 1'h0}; // @[PMDU.scala 1165:87]
  wire [30:0] _T_1375 = _T_1372[32] ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1376 = {_T_1375,_T_1372}; // @[Cat.scala 30:58]
  wire [63:0] _T_1377 = _T_476 ? _T_1371 : _T_1376; // @[PMDU.scala 1165:28]
  wire [63:0] _GEN_189 = _T_1354 == 16'h8000 & _T_1357 == 16'h8000 ? _T_1364 : _T_1377; // @[PMDU.scala 1161:70 1163:22 1165:22]
  wire [32:0] _T_1383 = {_GEN_189[31],_GEN_189[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1418 = io_out_bits_DecodeOut_ctrl_fuOpType[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1420 = _T_1418 ^ io_in_bits_Pctrl_mulres65_0[31:0]; // @[PMDU.scala 1187:74]
  wire [63:0] _T_1421 = io_out_bits_DecodeOut_ctrl_fuOpType[4] ? io_in_bits_Pctrl_mulres65_0[63:0] : {{32'd0}, _T_1420}; // @[PMDU.scala 1187:29]
  wire [70:0] _GEN_196 = io_in_bits_Pctrl_isC31 ? {{7'd0}, _T_1421} : _GEN_117; // @[PMDU.scala 1183:39 1187:23]
  wire [70:0] _GEN_201 = io_in_bits_Pctrl_isQ15orQ31 ? {{38'd0}, _T_1383} : _GEN_196; // @[PMDU.scala 1149:44 1168:23]
  wire [70:0] _GEN_205 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1289} : _GEN_201; // @[PMDU.scala 1126:40 1137:23]
  wire [70:0] _GEN_212 = io_in_bits_Pctrl_is3264 ? {{5'd0}, _T_1219} : _GEN_205; // @[PMDU.scala 1089:40 1099:23]
  wire [70:0] _GEN_230 = io_in_bits_Pctrl_is832 ? _GEN_117 : _GEN_212; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_236 = io_in_bits_Pctrl_isS1664 ? {{7'd0}, _T_1108} : _GEN_230; // @[PMDU.scala 1046:41 1048:19]
  wire [70:0] _GEN_263 = io_in_bits_Pctrl_isS1632 ? _GEN_117 : _GEN_236; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_280 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_117 : _GEN_263; // @[PMDU.scala 963:44]
  wire [70:0] adder68_1 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_117 : _GEN_280; // @[PMDU.scala 929:38]
  wire [70:0] _T_5 = adder68_0 + adder68_1; // @[PMDU.scala 726:24]
  wire  _T_949 = _T_538 & (_T_467 | _T_476) | _T_934; // @[PMDU.scala 1003:146]
  wire [33:0] _T_1045 = _T_949 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1031 = _T_929 ? 32'h0 : io_in_bits_Pctrl_mulres33_0[31:0]; // @[PMDU.scala 1016:102]
  wire [1:0] _T_1048 = _T_1031[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1049 = {_T_1048,_T_1031}; // @[Cat.scala 30:58]
  wire [33:0] _T_1050 = _T_1045 ^ _T_1049; // @[PMDU.scala 1022:56]
  wire [14:0] _T_1167 = io_in_bits_Pctrl_mulres17_1[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1168 = {_T_1167,io_in_bits_Pctrl_mulres17_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1169 = {15'h0,io_in_bits_Pctrl_mulres17_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_171 = _T_1156 ? _T_1168 : _T_1169; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_225 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_171} : 34'h0; // @[PMDU.scala 1051:39 1080:30]
  wire [33:0] _GEN_246 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_225; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_259 = io_in_bits_Pctrl_isS1632 ? _T_1050 : _GEN_246; // @[PMDU.scala 1000:41 1022:30]
  wire [33:0] _GEN_275 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_259; // @[PMDU.scala 963:44 981:30]
  wire [33:0] adder34_2_1 = io_in_bits_Pctrl_isMSW_3232 ? {{33'd0}, _T_687} : _GEN_275; // @[PMDU.scala 929:38 940:30]
  wire [31:0] _T_964 = _T_929 ? 32'h0 : io_in_bits_Pctrl_mulres17_0[31:0]; // @[PMDU.scala 1016:39]
  wire [1:0] _T_981 = _T_964[31] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_982 = {_T_981,_T_964}; // @[Cat.scala 30:58]
  wire [33:0] _T_983 = _T_1045 ^ _T_982; // @[PMDU.scala 1022:56]
  wire [14:0] _T_1128 = io_in_bits_Pctrl_mulres9_1[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1129 = {_T_1128,io_in_bits_Pctrl_mulres9_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1130 = {15'h0,io_in_bits_Pctrl_mulres9_1[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_167 = _T_1156 ? _T_1129 : _T_1130; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_220 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_167} : 34'h0; // @[PMDU.scala 1051:39 1080:30]
  wire [33:0] _GEN_241 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_220; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_254 = io_in_bits_Pctrl_isS1632 ? _T_983 : _GEN_241; // @[PMDU.scala 1000:41 1022:30]
  wire [33:0] _GEN_272 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_254; // @[PMDU.scala 963:44 981:30]
  wire [33:0] adder34_2_0 = io_in_bits_Pctrl_isMSW_3232 ? {{33'd0}, _T_687} : _GEN_272; // @[PMDU.scala 929:38 940:30]
  wire [70:0] _T_14 = {adder34_2_1,3'h0,adder34_2_0}; // @[Cat.scala 30:58]
  wire  _T_546 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h6 | _T_934; // @[PMDU.scala 906:59]
  wire [65:0] _T_567 = _T_546 ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_571 = io_in_bits_Pctrl_mulres65_0[63] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [65:0] _T_572 = {_T_571,io_in_bits_Pctrl_mulres65_0[63:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_573 = _T_567 ^ _T_572; // @[PMDU.scala 910:47]
  wire [70:0] _GEN_68 = io_in_bits_Pctrl_isPMA_64ONLY ? {{5'd0}, _T_573} : _T_14; // @[PMDU.scala 730:15 902:50 910:27]
  wire [70:0] _GEN_74 = io_in_bits_Pctrl_isQ63_64ONLY ? 71'h0 : _GEN_68; // @[PMDU.scala 886:50 890:27]
  wire [70:0] _GEN_81 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_14 : _GEN_74; // @[PMDU.scala 730:15 884:53]
  wire [70:0] _GEN_94 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_14 : _GEN_81; // @[PMDU.scala 730:15 836:50]
  wire [70:0] _GEN_106 = io_in_bits_Pctrl_isMul_8 ? _T_14 : _GEN_94; // @[PMDU.scala 730:15 779:45]
  wire [70:0] _GEN_118 = io_in_bits_Pctrl_isMul_16 ? _T_14 : _GEN_106; // @[PMDU.scala 730:15 735:40]
  wire [31:0] _T_1112 = io_in_bits_Pctrl_mulres33_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1113 = {_T_1112,io_in_bits_Pctrl_mulres33_0[31:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1209 = {io_in_bits_Pctrl_mulres65_0[64],io_in_bits_Pctrl_mulres65_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_1210 = {1'h0,io_in_bits_Pctrl_mulres65_0[64:0]}; // @[Cat.scala 30:58]
  wire [65:0] _GEN_175 = _T_1198 ? _T_1209 : _T_1210; // @[PMDU.scala 676:24 677:15 679:15]
  wire [65:0] _T_1222 = _T_1218 ^ _GEN_175; // @[PMDU.scala 1100:41]
  wire [31:0] _T_1274 = _T_467 ? 32'h0 : io_in_bits_Pctrl_mulres33_0[31:0]; // @[PMDU.scala 1134:23]
  wire [31:0] _T_1294 = _T_1274[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1295 = {_T_1294,_T_1274}; // @[Cat.scala 30:58]
  wire [63:0] _T_1296 = _T_1279 ^ _T_1295; // @[PMDU.scala 1138:50]
  wire [70:0] _GEN_197 = io_in_bits_Pctrl_isC31 ? {{70'd0}, io_out_bits_DecodeOut_ctrl_fuOpType[0]} : _GEN_118; // @[PMDU.scala 1183:39 1188:23]
  wire [70:0] _GEN_203 = io_in_bits_Pctrl_isQ15orQ31 ? _GEN_118 : _GEN_197; // @[PMDU.scala 1149:44]
  wire [70:0] _GEN_206 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1296} : _GEN_203; // @[PMDU.scala 1126:40 1138:23]
  wire [70:0] _GEN_213 = io_in_bits_Pctrl_is3264 ? {{5'd0}, _T_1222} : _GEN_206; // @[PMDU.scala 1089:40 1100:23]
  wire [70:0] _GEN_231 = io_in_bits_Pctrl_is832 ? _GEN_118 : _GEN_213; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_237 = io_in_bits_Pctrl_isS1664 ? {{7'd0}, _T_1113} : _GEN_231; // @[PMDU.scala 1046:41 1049:19]
  wire [70:0] _GEN_264 = io_in_bits_Pctrl_isS1632 ? _GEN_118 : _GEN_237; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_281 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_118 : _GEN_264; // @[PMDU.scala 963:44]
  wire [70:0] adder68_2 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_118 : _GEN_281; // @[PMDU.scala 929:38]
  wire [70:0] _T_7 = _T_5 + adder68_2; // @[PMDU.scala 726:36]
  wire [1:0] _T_1051 = _T_935 + _T_949; // @[PMDU.scala 1023:49]
  wire [14:0] _T_1174 = io_in_bits_Pctrl_mulres33_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1175 = {_T_1174,io_in_bits_Pctrl_mulres33_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1176 = {15'h0,io_in_bits_Pctrl_mulres33_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_172 = _T_1156 ? _T_1175 : _T_1176; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_226 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_172} : 34'h0; // @[PMDU.scala 1051:39 1081:30]
  wire [33:0] _GEN_247 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_226; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_260 = io_in_bits_Pctrl_isS1632 ? {{32'd0}, _T_1051} : _GEN_247; // @[PMDU.scala 1000:41 1023:30]
  wire [33:0] _GEN_278 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_260; // @[PMDU.scala 963:44]
  wire [33:0] adder34_3_1 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_278; // @[PMDU.scala 929:38]
  wire [14:0] _T_1135 = io_in_bits_Pctrl_mulres9_2[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1136 = {_T_1135,io_in_bits_Pctrl_mulres9_2[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1137 = {15'h0,io_in_bits_Pctrl_mulres9_2[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_168 = _T_1156 ? _T_1136 : _T_1137; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_221 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_168} : 34'h0; // @[PMDU.scala 1051:39 1081:30]
  wire [33:0] _GEN_242 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_221; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_255 = io_in_bits_Pctrl_isS1632 ? {{32'd0}, _T_1051} : _GEN_242; // @[PMDU.scala 1000:41 1023:30]
  wire [33:0] _GEN_277 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_255; // @[PMDU.scala 963:44]
  wire [33:0] adder34_3_0 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_277; // @[PMDU.scala 929:38]
  wire [70:0] _T_15 = {adder34_3_1,3'h0,adder34_3_0}; // @[Cat.scala 30:58]
  wire [1:0] _T_574 = _T_541 + _T_546; // @[PMDU.scala 911:46]
  wire [70:0] _GEN_69 = io_in_bits_Pctrl_isPMA_64ONLY ? {{69'd0}, _T_574} : _T_15; // @[PMDU.scala 731:15 902:50 911:27]
  wire [70:0] _GEN_77 = io_in_bits_Pctrl_isQ63_64ONLY ? _T_15 : _GEN_69; // @[PMDU.scala 731:15 886:50]
  wire [70:0] _GEN_83 = io_in_bits_Pctrl_isMul_32_64ONLY ? _T_15 : _GEN_77; // @[PMDU.scala 731:15 884:53]
  wire [70:0] _GEN_95 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_15 : _GEN_83; // @[PMDU.scala 731:15 836:50]
  wire [70:0] _GEN_107 = io_in_bits_Pctrl_isMul_8 ? _T_15 : _GEN_95; // @[PMDU.scala 731:15 779:45]
  wire [70:0] _GEN_119 = io_in_bits_Pctrl_isMul_16 ? _T_15 : _GEN_107; // @[PMDU.scala 731:15 735:40]
  wire [1:0] _T_1223 = {io_out_bits_DecodeOut_ctrl_fuOpType[0],1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1298 = _T_1266 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1272 = _T_467 ? io_in_bits_Pctrl_mulres65_0[31:0] : io_in_bits_Pctrl_mulres17_1[31:0]; // @[PMDU.scala 1133:23]
  wire [31:0] _T_1301 = _T_1272[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1302 = {_T_1301,_T_1272}; // @[Cat.scala 30:58]
  wire [63:0] _T_1303 = _T_1298 ^ _T_1302; // @[PMDU.scala 1139:50]
  wire [70:0] _GEN_207 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1303} : _GEN_119; // @[PMDU.scala 1126:40 1139:23]
  wire [70:0] _GEN_214 = io_in_bits_Pctrl_is3264 ? {{69'd0}, _T_1223} : _GEN_207; // @[PMDU.scala 1089:40 1101:23]
  wire [70:0] _GEN_232 = io_in_bits_Pctrl_is832 ? _GEN_119 : _GEN_214; // @[PMDU.scala 1051:39]
  wire [70:0] _GEN_249 = io_in_bits_Pctrl_isS1664 ? _GEN_119 : _GEN_232; // @[PMDU.scala 1046:41]
  wire [70:0] _GEN_267 = io_in_bits_Pctrl_isS1632 ? _GEN_119 : _GEN_249; // @[PMDU.scala 1000:41]
  wire [70:0] _GEN_284 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_119 : _GEN_267; // @[PMDU.scala 963:44]
  wire [70:0] adder68_3 = io_in_bits_Pctrl_isMSW_3232 ? _GEN_119 : _GEN_284; // @[PMDU.scala 929:38]
  wire [70:0] _T_9 = _T_7 + adder68_3; // @[PMDU.scala 726:48]
  wire [14:0] _T_1181 = io_in_bits_Pctrl_mulres65_0[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1182 = {_T_1181,io_in_bits_Pctrl_mulres65_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1183 = {15'h0,io_in_bits_Pctrl_mulres65_0[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_173 = _T_1156 ? _T_1182 : _T_1183; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_227 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_173} : 34'h0; // @[PMDU.scala 1051:39 1082:30]
  wire [33:0] _GEN_248 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_227; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_266 = io_in_bits_Pctrl_isS1632 ? 34'h0 : _GEN_248; // @[PMDU.scala 1000:41]
  wire [33:0] _GEN_283 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_266; // @[PMDU.scala 963:44]
  wire [33:0] adder34_4_1 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_283; // @[PMDU.scala 929:38]
  wire [14:0] _T_1142 = io_in_bits_Pctrl_mulres9_3[16] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1143 = {_T_1142,io_in_bits_Pctrl_mulres9_3[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_1144 = {15'h0,io_in_bits_Pctrl_mulres9_3[16:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_169 = _T_1156 ? _T_1143 : _T_1144; // @[PMDU.scala 676:24 677:15 679:15]
  wire [33:0] _GEN_222 = io_in_bits_Pctrl_is832 ? {{2'd0}, _GEN_169} : 34'h0; // @[PMDU.scala 1051:39 1082:30]
  wire [33:0] _GEN_243 = io_in_bits_Pctrl_isS1664 ? 34'h0 : _GEN_222; // @[PMDU.scala 1046:41]
  wire [33:0] _GEN_265 = io_in_bits_Pctrl_isS1632 ? 34'h0 : _GEN_243; // @[PMDU.scala 1000:41]
  wire [33:0] _GEN_282 = io_in_bits_Pctrl_isMSW_3216 ? 34'h0 : _GEN_265; // @[PMDU.scala 963:44]
  wire [33:0] adder34_4_0 = io_in_bits_Pctrl_isMSW_3232 ? 34'h0 : _GEN_282; // @[PMDU.scala 929:38]
  wire [70:0] _T_16 = {adder34_4_1,3'h0,adder34_4_0}; // @[Cat.scala 30:58]
  wire [31:0] _T_1276 = _T_467 ? 32'h0 : io_in_bits_Pctrl_mulres65_0[31:0]; // @[PMDU.scala 1135:23]
  wire [31:0] _T_1308 = _T_1276[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1309 = {_T_1308,_T_1276}; // @[Cat.scala 30:58]
  wire [63:0] _T_1310 = _T_1298 ^ _T_1309; // @[PMDU.scala 1140:50]
  wire [70:0] _GEN_208 = io_in_bits_Pctrl_is1664 ? {{7'd0}, _T_1310} : _T_16; // @[PMDU.scala 1126:40 1140:23 732:15]
  wire [70:0] _GEN_217 = io_in_bits_Pctrl_is3264 ? _T_16 : _GEN_208; // @[PMDU.scala 1089:40 732:15]
  wire [70:0] _GEN_234 = io_in_bits_Pctrl_is832 ? _T_16 : _GEN_217; // @[PMDU.scala 1051:39 732:15]
  wire [70:0] _GEN_251 = io_in_bits_Pctrl_isS1664 ? _T_16 : _GEN_234; // @[PMDU.scala 1046:41 732:15]
  wire [70:0] _GEN_268 = io_in_bits_Pctrl_isS1632 ? _T_16 : _GEN_251; // @[PMDU.scala 1000:41 732:15]
  wire [70:0] _GEN_285 = io_in_bits_Pctrl_isMSW_3216 ? _T_16 : _GEN_268; // @[PMDU.scala 732:15 963:44]
  wire [70:0] adder68_4 = io_in_bits_Pctrl_isMSW_3232 ? _T_16 : _GEN_285; // @[PMDU.scala 732:15 929:38]
  wire [70:0] tmp68 = _T_9 + adder68_4; // @[PMDU.scala 726:60]
  wire  _T_21 = io_out_bits_DecodeOut_ctrl_fuOpType[1:0] == 2'h1 | io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h9; // @[PMDU.scala 671:57]
  wire [15:0] _GEN_0 = _T_21 ? io_out_bits_DecodeOut_data_src2[31:16] : io_out_bits_DecodeOut_data_src2[15:0]; // @[PMDU.scala 687:23 689:29]
  wire [15:0] _GEN_1 = _T_21 ? io_out_bits_DecodeOut_data_src2[15:0] : io_out_bits_DecodeOut_data_src2[31:16]; // @[PMDU.scala 687:23 691:29]
  wire [15:0] _GEN_2 = _T_21 ? io_out_bits_DecodeOut_data_src2[63:48] : io_out_bits_DecodeOut_data_src2[47:32]; // @[PMDU.scala 687:23 689:29]
  wire [15:0] _GEN_3 = _T_21 ? io_out_bits_DecodeOut_data_src2[47:32] : io_out_bits_DecodeOut_data_src2[63:48]; // @[PMDU.scala 687:23 691:29]
  wire [63:0] _T_32 = {_GEN_3,_GEN_2,_GEN_1,_GEN_0}; // @[Cat.scala 30:58]
  wire  _T_34 = io_out_bits_DecodeOut_ctrl_fuOpType[1:0] == 2'h3; // @[PMDU.scala 672:44]
  wire [31:0] _T_48 = io_in_bits_Pctrl_mulres17_0[31:0]; // @[PMDU.scala 749:75]
  wire [16:0] _T_50 = _T_48[31:15]; // @[PMDU.scala 749:89]
  wire [31:0] _GEN_5 = _T_32[15:0] == 16'h8000 & io_out_bits_DecodeOut_data_src1[15:0] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_50}; // @[PMDU.scala 744:153 746:33 749:37]
  wire [31:0] _T_72 = io_in_bits_Pctrl_mulres17_1[31:0]; // @[PMDU.scala 751:75]
  wire [16:0] _T_74 = _T_72[31:15]; // @[PMDU.scala 751:89]
  wire [31:0] _GEN_7 = _T_32[31:16] == 16'h8000 & io_out_bits_DecodeOut_data_src1[31:16] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_74}; // @[PMDU.scala 744:153 746:33 751:37]
  wire [31:0] _T_96 = io_in_bits_Pctrl_mulres33_0[31:0]; // @[PMDU.scala 753:75]
  wire [16:0] _T_98 = _T_96[31:15]; // @[PMDU.scala 753:89]
  wire [31:0] _GEN_9 = _T_32[47:32] == 16'h8000 & io_out_bits_DecodeOut_data_src1[47:32] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_98}; // @[PMDU.scala 744:153 746:33 753:37]
  wire  _GEN_10 = _T_32[63:48] == 16'h8000 & io_out_bits_DecodeOut_data_src1[63:48] == 16'h8000 | (_T_32[47:32] == 16'h8000
     & io_out_bits_DecodeOut_data_src1[47:32] == 16'h8000 | (_T_32[31:16] == 16'h8000 & io_out_bits_DecodeOut_data_src1[
    31:16] == 16'h8000 | _T_32[15:0] == 16'h8000 & io_out_bits_DecodeOut_data_src1[15:0] == 16'h8000)); // @[PMDU.scala 744:153 745:59]
  wire [31:0] _GEN_11 = _T_32[63:48] == 16'h8000 & io_out_bits_DecodeOut_data_src1[63:48] == 16'h8000 ? 32'h7fff : {{15
    'd0}, _T_1367}; // @[PMDU.scala 744:153 746:33 755:37]
  wire [63:0] _T_133 = {_GEN_11[15:0],_GEN_9[15:0],_GEN_7[15:0],_GEN_5[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_136 = {io_in_bits_Pctrl_mulres65_0[31:0],io_in_bits_Pctrl_mulres17_0[31:0]}; // @[Cat.scala 30:58]
  wire  _GEN_12 = _T_34 & _GEN_10; // @[PMDU.scala 705:35 738:39]
  wire [63:0] _GEN_13 = _T_34 ? _T_133 : _T_136; // @[PMDU.scala 738:39 739:36 764:36]
  wire [7:0] _GEN_14 = _T_21 ? io_out_bits_DecodeOut_data_src2[15:8] : io_out_bits_DecodeOut_data_src2[7:0]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_15 = _T_21 ? io_out_bits_DecodeOut_data_src2[7:0] : io_out_bits_DecodeOut_data_src2[15:8]; // @[PMDU.scala 687:23 691:29]
  wire [7:0] _GEN_16 = _T_21 ? io_out_bits_DecodeOut_data_src2[31:24] : io_out_bits_DecodeOut_data_src2[23:16]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_17 = _T_21 ? io_out_bits_DecodeOut_data_src2[23:16] : io_out_bits_DecodeOut_data_src2[31:24]; // @[PMDU.scala 687:23 691:29]
  wire [7:0] _GEN_18 = _T_21 ? io_out_bits_DecodeOut_data_src2[47:40] : io_out_bits_DecodeOut_data_src2[39:32]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_19 = _T_21 ? io_out_bits_DecodeOut_data_src2[39:32] : io_out_bits_DecodeOut_data_src2[47:40]; // @[PMDU.scala 687:23 691:29]
  wire [7:0] _GEN_20 = _T_21 ? io_out_bits_DecodeOut_data_src2[63:56] : io_out_bits_DecodeOut_data_src2[55:48]; // @[PMDU.scala 687:23 689:29]
  wire [7:0] _GEN_21 = _T_21 ? io_out_bits_DecodeOut_data_src2[55:48] : io_out_bits_DecodeOut_data_src2[63:56]; // @[PMDU.scala 687:23 691:29]
  wire [63:0] _T_164 = {_GEN_21,_GEN_20,_GEN_19,_GEN_18,_GEN_17,_GEN_16,_GEN_15,_GEN_14}; // @[Cat.scala 30:58]
  wire [15:0] _T_180 = io_in_bits_Pctrl_mulres9_0[15:0]; // @[PMDU.scala 793:74]
  wire [8:0] _T_182 = _T_180[15:7]; // @[PMDU.scala 793:87]
  wire [15:0] _GEN_23 = _T_164[7:0] == 8'h80 & io_out_bits_DecodeOut_data_src1[7:0] == 8'h80 ? 16'h7f : {{7'd0}, _T_182}
    ; // @[PMDU.scala 788:151 790:33 793:37]
  wire [15:0] _T_204 = io_in_bits_Pctrl_mulres9_1[15:0]; // @[PMDU.scala 795:74]
  wire [8:0] _T_206 = _T_204[15:7]; // @[PMDU.scala 795:87]
  wire [15:0] _GEN_25 = _T_164[15:8] == 8'h80 & io_out_bits_DecodeOut_data_src1[15:8] == 8'h80 ? 16'h7f : {{7'd0},
    _T_206}; // @[PMDU.scala 788:151 790:33 795:37]
  wire [15:0] _T_228 = io_in_bits_Pctrl_mulres9_2[15:0]; // @[PMDU.scala 797:74]
  wire [8:0] _T_230 = _T_228[15:7]; // @[PMDU.scala 797:87]
  wire [15:0] _GEN_27 = _T_164[23:16] == 8'h80 & io_out_bits_DecodeOut_data_src1[23:16] == 8'h80 ? 16'h7f : {{7'd0},
    _T_230}; // @[PMDU.scala 788:151 790:33 797:37]
  wire [15:0] _T_252 = io_in_bits_Pctrl_mulres9_3[15:0]; // @[PMDU.scala 799:74]
  wire [8:0] _T_254 = _T_252[15:7]; // @[PMDU.scala 799:87]
  wire [15:0] _GEN_29 = _T_164[31:24] == 8'h80 & io_out_bits_DecodeOut_data_src1[31:24] == 8'h80 ? 16'h7f : {{7'd0},
    _T_254}; // @[PMDU.scala 788:151 790:33 799:37]
  wire [15:0] _T_276 = io_in_bits_Pctrl_mulres17_0[15:0]; // @[PMDU.scala 801:75]
  wire [8:0] _T_278 = _T_276[15:7]; // @[PMDU.scala 801:88]
  wire [15:0] _GEN_31 = _T_164[39:32] == 8'h80 & io_out_bits_DecodeOut_data_src1[39:32] == 8'h80 ? 16'h7f : {{7'd0},
    _T_278}; // @[PMDU.scala 788:151 790:33 801:37]
  wire [15:0] _T_300 = io_in_bits_Pctrl_mulres17_1[15:0]; // @[PMDU.scala 803:75]
  wire [8:0] _T_302 = _T_300[15:7]; // @[PMDU.scala 803:88]
  wire [15:0] _GEN_33 = _T_164[47:40] == 8'h80 & io_out_bits_DecodeOut_data_src1[47:40] == 8'h80 ? 16'h7f : {{7'd0},
    _T_302}; // @[PMDU.scala 788:151 790:33 803:37]
  wire [15:0] _T_324 = io_in_bits_Pctrl_mulres33_0[15:0]; // @[PMDU.scala 805:75]
  wire [8:0] _T_326 = _T_324[15:7]; // @[PMDU.scala 805:88]
  wire  _GEN_34 = _T_164[55:48] == 8'h80 & io_out_bits_DecodeOut_data_src1[55:48] == 8'h80 | (_T_164[47:40] == 8'h80 &
    io_out_bits_DecodeOut_data_src1[47:40] == 8'h80 | (_T_164[39:32] == 8'h80 & io_out_bits_DecodeOut_data_src1[39:32]
     == 8'h80 | (_T_164[31:24] == 8'h80 & io_out_bits_DecodeOut_data_src1[31:24] == 8'h80 | (_T_164[23:16] == 8'h80 &
    io_out_bits_DecodeOut_data_src1[23:16] == 8'h80 | (_T_164[15:8] == 8'h80 & io_out_bits_DecodeOut_data_src1[15:8] == 8'h80
     | _T_164[7:0] == 8'h80 & io_out_bits_DecodeOut_data_src1[7:0] == 8'h80))))); // @[PMDU.scala 788:151 789:59]
  wire [15:0] _GEN_35 = _T_164[55:48] == 8'h80 & io_out_bits_DecodeOut_data_src1[55:48] == 8'h80 ? 16'h7f : {{7'd0},
    _T_326}; // @[PMDU.scala 788:151 790:33 805:37]
  wire [15:0] _T_348 = io_in_bits_Pctrl_mulres65_0[15:0]; // @[PMDU.scala 807:75]
  wire [8:0] _T_350 = _T_348[15:7]; // @[PMDU.scala 807:88]
  wire  _GEN_36 = _T_164[63:56] == 8'h80 & io_out_bits_DecodeOut_data_src1[63:56] == 8'h80 | _GEN_34; // @[PMDU.scala 788:151 789:59]
  wire [15:0] _GEN_37 = _T_164[63:56] == 8'h80 & io_out_bits_DecodeOut_data_src1[63:56] == 8'h80 ? 16'h7f : {{7'd0},
    _T_350}; // @[PMDU.scala 788:151 790:33 807:37]
  wire [63:0] _T_365 = {_GEN_37[7:0],_GEN_35[7:0],_GEN_33[7:0],_GEN_31[7:0],_GEN_29[7:0],_GEN_27[7:0],_GEN_25[7:0],
    _GEN_23[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_400 = {io_in_bits_Pctrl_mulres65_0[15:0],io_in_bits_Pctrl_mulres9_2[15:0],io_in_bits_Pctrl_mulres9_1[15
    :0],io_in_bits_Pctrl_mulres9_0[15:0]}; // @[Cat.scala 30:58]
  wire  _GEN_38 = _T_34 & _GEN_36; // @[PMDU.scala 705:35 782:39]
  wire [63:0] _GEN_39 = _T_34 ? _T_365 : _T_400; // @[PMDU.scala 782:39 783:36 816:36]
  wire [32:0] _T_445 = tmp68[32] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _GEN_304 = {{1'd0}, _T_445}; // @[PMDU.scala 870:63]
  wire [33:0] _T_447 = _GEN_304 ^ tmp68[33:0]; // @[PMDU.scala 870:63]
  wire  _T_449 = _T_447[32:31] != 2'h0; // @[PMDU.scala 870:92]
  wire [31:0] _GEN_44 = tmp68[32] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 872:65 873:36 875:37]
  wire  _GEN_45 = _T_447[32:31] != 2'h0 | _T_422; // @[PMDU.scala 870:100 871:59]
  wire [31:0] _GEN_46 = _T_447[32:31] != 2'h0 ? _GEN_44 : tmp68[31:0]; // @[PMDU.scala 870:100]
  wire  _GEN_47 = _T_467 ? _GEN_45 : _T_422; // @[PMDU.scala 869:53]
  wire [31:0] _GEN_48 = _T_467 ? _GEN_46 : tmp68[31:0]; // @[PMDU.scala 869:53]
  wire  _GEN_51 = _T_461 == 16'h8000 & _T_464 == 16'h8000 | _GEN_47; // @[PMDU.scala 851:77 852:55]
  wire [32:0] _T_497 = tmp68[69] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _GEN_305 = {{1'd0}, _T_497}; // @[PMDU.scala 870:63]
  wire [33:0] _T_499 = _GEN_305 ^ tmp68[70:37]; // @[PMDU.scala 870:63]
  wire  _T_501 = _T_499[32:31] != 2'h0; // @[PMDU.scala 870:92]
  wire [31:0] _GEN_53 = tmp68[69] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 872:65 873:36 875:37]
  wire  _GEN_54 = _T_499[32:31] != 2'h0 | _GEN_51; // @[PMDU.scala 870:100 871:59]
  wire [31:0] _GEN_55 = _T_499[32:31] != 2'h0 ? _GEN_53 : tmp68[68:37]; // @[PMDU.scala 870:100]
  wire  _GEN_56 = _T_467 ? _GEN_54 : _GEN_51; // @[PMDU.scala 869:53]
  wire [31:0] _GEN_57 = _T_467 ? _GEN_55 : tmp68[68:37]; // @[PMDU.scala 869:53]
  wire [63:0] _T_509 = {_GEN_57,_GEN_48}; // @[Cat.scala 30:58]
  wire [64:0] _T_519 = tmp68[64] ? 65'h1ffffffffffffffff : 65'h0; // @[Bitwise.scala 72:12]
  wire [70:0] _GEN_306 = {{6'd0}, _T_519}; // @[PMDU.scala 892:41]
  wire [70:0] _T_520 = _GEN_306 ^ tmp68; // @[PMDU.scala 892:41]
  wire  _T_522 = _T_520[64:63] != 2'h0; // @[PMDU.scala 892:56]
  wire [63:0] _GEN_58 = tmp68[64] ? 64'h8000000000000000 : 64'h7fffffffffffffff; // @[PMDU.scala 894:43 895:29 897:29]
  wire [63:0] _GEN_60 = _T_520[64:63] != 2'h0 ? _GEN_58 : tmp68[63:0]; // @[PMDU.scala 892:64]
  wire  _T_552 = ~(_T_924 & _T_467); // @[PMDU.scala 907:34]
  wire [65:0] _T_578 = tmp68[65] ? 66'h3ffffffffffffffff : 66'h0; // @[Bitwise.scala 72:12]
  wire [70:0] _GEN_307 = {{5'd0}, _T_578}; // @[PMDU.scala 914:45]
  wire [70:0] _T_579 = _GEN_307 ^ tmp68; // @[PMDU.scala 914:45]
  wire  _T_581 = _T_579[65:63] != 3'h0; // @[PMDU.scala 914:59]
  wire [63:0] _GEN_61 = tmp68[65] ? 64'h8000000000000000 : 64'h7fffffffffffffff; // @[PMDU.scala 916:40 917:33 919:33]
  wire [63:0] _GEN_63 = _T_579[65:63] != 3'h0 ? _GEN_61 : tmp68[63:0]; // @[PMDU.scala 914:66]
  wire  _GEN_64 = _T_552 & _T_581; // @[PMDU.scala 913:33 705:35]
  wire [63:0] _GEN_65 = _T_552 ? _GEN_63 : tmp68[63:0]; // @[PMDU.scala 913:33]
  wire  _GEN_70 = io_in_bits_Pctrl_isPMA_64ONLY & _GEN_64; // @[PMDU.scala 705:35 902:50]
  wire [63:0] _GEN_71 = io_in_bits_Pctrl_isPMA_64ONLY ? _GEN_65 : 64'h0; // @[PMDU.scala 704:24 902:50 903:32]
  wire  _GEN_75 = io_in_bits_Pctrl_isQ63_64ONLY ? _T_522 : _GEN_70; // @[PMDU.scala 886:50]
  wire [63:0] _GEN_76 = io_in_bits_Pctrl_isQ63_64ONLY ? _GEN_60 : _GEN_71; // @[PMDU.scala 886:50 887:32]
  wire [63:0] _GEN_78 = io_in_bits_Pctrl_isMul_32_64ONLY ? io_in_bits_Pctrl_mulres65_0[63:0] : _GEN_76; // @[PMDU.scala 884:53 885:32]
  wire  _GEN_82 = io_in_bits_Pctrl_isMul_32_64ONLY ? 1'h0 : _GEN_75; // @[PMDU.scala 705:35 884:53]
  wire  _GEN_84 = io_in_bits_Pctrl_isQ15_64ONLY ? _GEN_56 : _GEN_82; // @[PMDU.scala 836:50]
  wire [63:0] _GEN_91 = io_in_bits_Pctrl_isQ15_64ONLY ? _T_509 : _GEN_78; // @[PMDU.scala 836:50 837:32]
  wire  _GEN_96 = io_in_bits_Pctrl_isMul_8 ? _GEN_38 : _GEN_84; // @[PMDU.scala 779:45]
  wire [63:0] _GEN_97 = io_in_bits_Pctrl_isMul_8 ? _GEN_39 : _GEN_91; // @[PMDU.scala 779:45]
  wire  _GEN_108 = io_in_bits_Pctrl_isMul_16 ? _GEN_12 : _GEN_96; // @[PMDU.scala 735:40]
  wire [63:0] _GEN_109 = io_in_bits_Pctrl_isMul_16 ? _GEN_13 : _GEN_97; // @[PMDU.scala 735:40]
  wire  _T_612 = _T_694 & io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h0; // @[PMDU.scala 934:52]
  wire  _GEN_121 = _T_449 | _GEN_108; // @[PMDU.scala 945:96 946:55]
  wire  _GEN_123 = _T_803 & io_out_bits_DecodeOut_data_src2[31:0] == 32'h80000000 | _GEN_108; // @[PMDU.scala 954:147 955:55]
  wire [31:0] _GEN_124 = _T_803 & io_out_bits_DecodeOut_data_src2[31:0] == 32'h80000000 ? 32'h7fffffff : tmp68[31:0]; // @[PMDU.scala 954:147 956:29]
  wire  _GEN_125 = _T_697 ? _GEN_123 : _GEN_108; // @[PMDU.scala 953:32]
  wire [31:0] _GEN_126 = _T_697 ? _GEN_124 : tmp68[31:0]; // @[PMDU.scala 953:32]
  wire  _GEN_127 = _T_612 | _T_687 ? _GEN_121 : _GEN_125; // @[PMDU.scala 944:33]
  wire [31:0] _GEN_128 = _T_612 | _T_687 ? _GEN_46 : _GEN_126; // @[PMDU.scala 944:33]
  wire  _GEN_130 = _T_501 | _GEN_127; // @[PMDU.scala 945:96 946:55]
  wire  _GEN_132 = _T_880 & io_out_bits_DecodeOut_data_src2[63:32] == 32'h80000000 | _GEN_127; // @[PMDU.scala 954:147 955:55]
  wire [31:0] _GEN_133 = _T_880 & io_out_bits_DecodeOut_data_src2[63:32] == 32'h80000000 ? 32'h7fffffff : tmp68[68:37]; // @[PMDU.scala 954:147 956:29]
  wire  _GEN_134 = _T_697 ? _GEN_132 : _GEN_127; // @[PMDU.scala 953:32]
  wire [31:0] _GEN_135 = _T_697 ? _GEN_133 : tmp68[68:37]; // @[PMDU.scala 953:32]
  wire  _GEN_136 = _T_612 | _T_687 ? _GEN_130 : _GEN_134; // @[PMDU.scala 944:33]
  wire [31:0] _GEN_137 = _T_612 | _T_687 ? _GEN_55 : _GEN_135; // @[PMDU.scala 944:33]
  wire [63:0] _T_763 = {_GEN_137,_GEN_128}; // @[Cat.scala 30:58]
  wire  _T_768 = io_out_bits_DecodeOut_ctrl_fuOpType[2:0] == 3'h3 | io_out_bits_DecodeOut_ctrl_fuOpType[6:5] == 2'h3; // @[PMDU.scala 967:54]
  wire  _GEN_138 = _T_847 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80000000 & _T_781 == 16'h8000 | _GEN_108; // @[PMDU.scala 975:127 976:51]
  wire  _GEN_141 = _T_449 | _GEN_138; // @[PMDU.scala 987:96 988:55]
  wire  _GEN_143 = _T_768 ? _GEN_141 : _GEN_138; // @[PMDU.scala 986:26]
  wire [31:0] _GEN_144 = _T_768 ? _GEN_46 : tmp68[31:0]; // @[PMDU.scala 986:26]
  wire  _GEN_145 = _T_847 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80000000 & _T_858 == 16'h8000 | _GEN_143; // @[PMDU.scala 975:127 976:51]
  wire  _GEN_148 = _T_501 | _GEN_145; // @[PMDU.scala 987:96 988:55]
  wire  _GEN_150 = _T_768 ? _GEN_148 : _GEN_145; // @[PMDU.scala 986:26]
  wire [31:0] _GEN_151 = _T_768 ? _GEN_55 : tmp68[68:37]; // @[PMDU.scala 986:26]
  wire [63:0] _T_918 = {_GEN_151,_GEN_144}; // @[Cat.scala 30:58]
  wire  _T_951 = io_out_bits_DecodeOut_ctrl_fuOpType[6:1] == 6'he; // @[PMDU.scala 1004:40]
  wire  _T_959 = io_out_bits_DecodeOut_ctrl_fuOpType[6:3] == 4'h4 | _T_922 | _T_476; // @[PMDU.scala 1005:84]
  wire [31:0] _GEN_152 = _T_951 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80008000 &
    io_out_bits_DecodeOut_data_src2[31:0] == 32'h80008000 ? 32'h7fffffff : tmp68[31:0]; // @[PMDU.scala 1025:21 1026:211 1027:25]
  wire  _GEN_153 = _T_951 & io_out_bits_DecodeOut_data_src1[31:0] == 32'h80008000 & io_out_bits_DecodeOut_data_src2[31:0
    ] == 32'h80008000 | _GEN_108; // @[PMDU.scala 1026:211 1028:51]
  wire [33:0] _T_1008 = tmp68[33] ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1010 = _T_1008 ^ tmp68[33:0]; // @[PMDU.scala 1031:59]
  wire [31:0] _GEN_154 = tmp68[33] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 1033:61 1034:33 1036:33]
  wire  _GEN_155 = _T_1010[33:31] != 3'h0 | _GEN_153; // @[PMDU.scala 1031:96 1032:55]
  wire [31:0] _GEN_156 = _T_1010[33:31] != 3'h0 ? _GEN_154 : _GEN_152; // @[PMDU.scala 1031:96]
  wire  _GEN_157 = _T_959 ? _GEN_155 : _GEN_153; // @[PMDU.scala 1030:33]
  wire [31:0] _GEN_158 = _T_959 ? _GEN_156 : _GEN_152; // @[PMDU.scala 1030:33]
  wire [31:0] _GEN_159 = _T_951 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80008000 &
    io_out_bits_DecodeOut_data_src2[63:32] == 32'h80008000 ? 32'h7fffffff : tmp68[68:37]; // @[PMDU.scala 1025:21 1026:211 1027:25]
  wire  _GEN_160 = _T_951 & io_out_bits_DecodeOut_data_src1[63:32] == 32'h80008000 & io_out_bits_DecodeOut_data_src2[63:
    32] == 32'h80008000 | _GEN_157; // @[PMDU.scala 1026:211 1028:51]
  wire [33:0] _T_1075 = tmp68[70] ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12]
  wire [33:0] _T_1077 = _T_1075 ^ tmp68[70:37]; // @[PMDU.scala 1031:59]
  wire [31:0] _GEN_161 = tmp68[70] ? 32'h80000000 : 32'h7fffffff; // @[PMDU.scala 1033:61 1034:33 1036:33]
  wire  _GEN_162 = _T_1077[33:31] != 3'h0 | _GEN_160; // @[PMDU.scala 1031:96 1032:55]
  wire [31:0] _GEN_163 = _T_1077[33:31] != 3'h0 ? _GEN_161 : _GEN_159; // @[PMDU.scala 1031:96]
  wire  _GEN_164 = _T_959 ? _GEN_162 : _GEN_160; // @[PMDU.scala 1030:33]
  wire [31:0] _GEN_165 = _T_959 ? _GEN_163 : _GEN_159; // @[PMDU.scala 1030:33]
  wire [63:0] _T_1096 = {_GEN_165,_GEN_158}; // @[Cat.scala 30:58]
  wire [63:0] _T_1195 = {tmp68[68:37],tmp68[31:0]}; // @[Cat.scala 30:58]
  wire  _GEN_178 = _T_581 | _GEN_108; // @[PMDU.scala 1105:68 1106:55]
  wire  _GEN_180 = ~io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65:64] != 2'h0 | _GEN_108; // @[PMDU.scala 1117:61 1118:55]
  wire [63:0] _GEN_181 = ~io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65:64] != 2'h0 ? 64'hffffffffffffffff : tmp68[
    63:0]; // @[PMDU.scala 1117:61 1119:29]
  wire  _GEN_182 = io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65] | _GEN_180; // @[PMDU.scala 1114:52 1115:55]
  wire [63:0] _GEN_183 = io_out_bits_DecodeOut_ctrl_fuOpType[0] & tmp68[65] ? 64'h0 : _GEN_181; // @[PMDU.scala 1114:52 1116:29]
  wire  _GEN_184 = _T_1198 ? _GEN_178 : _GEN_182; // @[PMDU.scala 1104:31]
  wire [63:0] _GEN_185 = _T_1198 ? _GEN_63 : _GEN_183; // @[PMDU.scala 1104:31]
  wire  _GEN_186 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _GEN_184 : _GEN_108; // @[PMDU.scala 1103:29]
  wire [63:0] _GEN_187 = io_out_bits_DecodeOut_ctrl_fuOpType[3] ? _GEN_185 : tmp68[63:0]; // @[PMDU.scala 1103:29]
  wire  _GEN_188 = _T_1354 == 16'h8000 & _T_1357 == 16'h8000 | _GEN_108; // @[PMDU.scala 1161:70 1162:47]
  wire [31:0] _T_1387 = tmp68[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1388 = {_T_1387,tmp68[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1391 = tmp68[32] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [70:0] _GEN_313 = {{38'd0}, _T_1391}; // @[PMDU.scala 1172:41]
  wire [70:0] _T_1392 = _GEN_313 ^ tmp68; // @[PMDU.scala 1172:41]
  wire [63:0] _GEN_190 = tmp68[32] ? 64'hffffffff80000000 : 64'h7fffffff; // @[PMDU.scala 1174:43 1175:29 1177:29]
  wire  _GEN_191 = _T_1392[32:31] != 2'h0 | _GEN_188; // @[PMDU.scala 1172:64 1173:51]
  wire [63:0] _GEN_192 = _T_1392[32:31] != 2'h0 ? _GEN_190 : _T_1388; // @[PMDU.scala 1171:21 1172:64]
  wire [63:0] _GEN_193 = _T_686 ? _GEN_192 : _GEN_189; // @[PMDU.scala 1170:30]
  wire  _GEN_194 = _T_686 ? _GEN_191 : _GEN_188; // @[PMDU.scala 1170:30]
  wire [63:0] _T_1431 = io_out_bits_DecodeOut_ctrl_fuOpType[4] ? tmp68[63:0] : _T_1388; // @[PMDU.scala 1189:16]
  wire [63:0] _GEN_198 = io_in_bits_Pctrl_isC31 ? _T_1431 : _GEN_109; // @[PMDU.scala 1183:39 1184:28]
  wire  _GEN_199 = io_in_bits_Pctrl_isQ15orQ31 ? _GEN_194 : _GEN_108; // @[PMDU.scala 1149:44]
  wire [63:0] _GEN_202 = io_in_bits_Pctrl_isQ15orQ31 ? _GEN_193 : _GEN_198; // @[PMDU.scala 1149:44 1150:28]
  wire [63:0] _GEN_209 = io_in_bits_Pctrl_is1664 ? tmp68[63:0] : _GEN_202; // @[PMDU.scala 1126:40 1130:28]
  wire  _GEN_210 = io_in_bits_Pctrl_is1664 ? _GEN_108 : _GEN_199; // @[PMDU.scala 1126:40]
  wire  _GEN_215 = io_in_bits_Pctrl_is3264 ? _GEN_186 : _GEN_210; // @[PMDU.scala 1089:40]
  wire [63:0] _GEN_216 = io_in_bits_Pctrl_is3264 ? _GEN_187 : _GEN_209; // @[PMDU.scala 1089:40 1093:28]
  wire [63:0] _GEN_228 = io_in_bits_Pctrl_is832 ? _T_1195 : _GEN_216; // @[PMDU.scala 1051:39 1053:28]
  wire  _GEN_233 = io_in_bits_Pctrl_is832 ? _GEN_108 : _GEN_215; // @[PMDU.scala 1051:39]
  wire [63:0] _GEN_238 = io_in_bits_Pctrl_isS1664 ? tmp68[63:0] : _GEN_228; // @[PMDU.scala 1046:41 1050:28]
  wire  _GEN_250 = io_in_bits_Pctrl_isS1664 ? _GEN_108 : _GEN_233; // @[PMDU.scala 1046:41]
  wire  _GEN_256 = io_in_bits_Pctrl_isS1632 ? _GEN_164 : _GEN_250; // @[PMDU.scala 1000:41]
  wire [63:0] _GEN_261 = io_in_bits_Pctrl_isS1632 ? _T_1096 : _GEN_238; // @[PMDU.scala 1000:41 1006:28]
  wire  _GEN_269 = io_in_bits_Pctrl_isMSW_3216 ? _GEN_150 : _GEN_256; // @[PMDU.scala 963:44]
  wire [63:0] _GEN_276 = io_in_bits_Pctrl_isMSW_3216 ? _T_918 : _GEN_261; // @[PMDU.scala 963:44 964:28]
  assign io_in_ready = _T | ~io_in_valid; // @[PMDU.scala 701:35]
  assign io_out_valid = io_in_valid; // @[PMDU.scala 700:18]
  assign io_out_bits_result = io_in_bits_Pctrl_isMSW_3232 ? _T_763 : _GEN_276; // @[PMDU.scala 929:38 930:28]
  assign io_out_bits_DecodeOut_cf_pc = io_in_bits_DecodeIn_cf_pc; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_cf_runahead_checkpoint_id = io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_ctrl_fuOpType = io_in_bits_DecodeIn_ctrl_fuOpType; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_ctrl_rfWen = io_in_bits_DecodeIn_ctrl_rfWen; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_ctrl_rfDest = io_in_bits_DecodeIn_ctrl_rfDest; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_data_src1 = io_in_bits_DecodeIn_data_src1; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_data_src2 = io_in_bits_DecodeIn_data_src2; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_data_src3 = io_in_bits_DecodeIn_data_src3; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_pext_OV = io_in_bits_Pctrl_isMSW_3232 ? _GEN_136 : _GEN_269; // @[PMDU.scala 929:38]
  assign io_out_bits_DecodeOut_InstNo = io_in_bits_DecodeIn_InstNo; // @[PMDU.scala 703:27]
  assign io_out_bits_DecodeOut_InstFlag = io_in_bits_DecodeIn_InstFlag; // @[PMDU.scala 703:27]
  assign io_FirstStageFire = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
endmodule
module MulAdd_onestage(
  input  [16:0] io_in_srcs_0,
  input  [16:0] io_in_srcs_1,
  output [33:0] io_out_result
);
  assign io_out_result = $signed(io_in_srcs_0) * $signed(io_in_srcs_1); // @[PIDU.scala 138:44]
endmodule
module MulAdd_onestage_2(
  input  [32:0] io_in_srcs_0,
  input  [32:0] io_in_srcs_1,
  output [65:0] io_out_result
);
  assign io_out_result = $signed(io_in_srcs_0) * $signed(io_in_srcs_1); // @[PIDU.scala 138:44]
endmodule
module MulAdd_onestage_3(
  input  [64:0]  io_in_srcs_0,
  input  [64:0]  io_in_srcs_1,
  output [129:0] io_out_result
);
  assign io_out_result = $signed(io_in_srcs_0) * $signed(io_in_srcs_1); // @[PIDU.scala 138:44]
endmodule
module MulAdd_onestage_4(
  input  [8:0]  io_in_srcs_0,
  input  [8:0]  io_in_srcs_1,
  output [17:0] io_out_result
);
  assign io_out_result = $signed(io_in_srcs_0) * $signed(io_in_srcs_1); // @[PIDU.scala 138:44]
endmodule
module PIDU(
  input  [63:0]  io_DecodeIn_cf_instr,
  input  [4:0]   io_DecodeIn_cf_instrType,
  input  [6:0]   io_DecodeIn_ctrl_fuOpType,
  input  [2:0]   io_DecodeIn_ctrl_funct3,
  input          io_DecodeIn_ctrl_func24,
  input          io_DecodeIn_ctrl_func23,
  input  [63:0]  io_DecodeIn_data_src1,
  input  [63:0]  io_DecodeIn_data_src2,
  output         io_Pctrl_isAdd_64,
  output         io_Pctrl_isAdd_32,
  output         io_Pctrl_isAdd_16,
  output         io_Pctrl_isAdd_8,
  output         io_Pctrl_isAdd_Q15,
  output         io_Pctrl_isAdd_Q31,
  output         io_Pctrl_isAdd_C31,
  output         io_Pctrl_isAve,
  output         io_Pctrl_isAdd,
  output         io_Pctrl_isSub_64,
  output         io_Pctrl_isSub_32,
  output         io_Pctrl_isSub_16,
  output         io_Pctrl_isSub_8,
  output         io_Pctrl_isSub_Q15,
  output         io_Pctrl_isSub_Q31,
  output         io_Pctrl_isSub_C31,
  output         io_Pctrl_isCras_16,
  output         io_Pctrl_isCrsa_16,
  output         io_Pctrl_isCras_32,
  output         io_Pctrl_isCrsa_32,
  output         io_Pctrl_isCr,
  output         io_Pctrl_isStas_16,
  output         io_Pctrl_isStsa_16,
  output         io_Pctrl_isStas_32,
  output         io_Pctrl_isStsa_32,
  output         io_Pctrl_isSt,
  output         io_Pctrl_isComp_16,
  output         io_Pctrl_isComp_8,
  output         io_Pctrl_isCompare,
  output         io_Pctrl_isMaxMin_16,
  output         io_Pctrl_isMaxMin_8,
  output         io_Pctrl_isMaxMin_XLEN,
  output         io_Pctrl_isMaxMin_32,
  output         io_Pctrl_isMaxMin,
  output         io_Pctrl_isPbs,
  output         io_Pctrl_isRs_16,
  output         io_Pctrl_isLs_16,
  output         io_Pctrl_isLR_16,
  output         io_Pctrl_isRs_8,
  output         io_Pctrl_isLs_8,
  output         io_Pctrl_isLR_8,
  output         io_Pctrl_isRs_32,
  output         io_Pctrl_isLs_32,
  output         io_Pctrl_isLR_32,
  output         io_Pctrl_isLR_Q31,
  output         io_Pctrl_isLs_Q31,
  output         io_Pctrl_isRs_XLEN,
  output         io_Pctrl_isSRAIWU,
  output         io_Pctrl_isFSRW,
  output         io_Pctrl_isWext,
  output         io_Pctrl_isShifter,
  output         io_Pctrl_isClip_16,
  output         io_Pctrl_isClip_8,
  output         io_Pctrl_isclip_32,
  output         io_Pctrl_isClip,
  output         io_Pctrl_isSat_16,
  output         io_Pctrl_isSat_8,
  output         io_Pctrl_isSat_32,
  output         io_Pctrl_isSat_W,
  output         io_Pctrl_isSat,
  output         io_Pctrl_isCnt_16,
  output         io_Pctrl_isCnt_8,
  output         io_Pctrl_isCnt_32,
  output         io_Pctrl_isCnt,
  output         io_Pctrl_isSwap_16,
  output         io_Pctrl_isSwap_8,
  output         io_Pctrl_isSwap,
  output         io_Pctrl_isUnpack,
  output         io_Pctrl_isBitrev,
  output         io_Pctrl_isCmix,
  output         io_Pctrl_isInsertb,
  output         io_Pctrl_isPackbb,
  output         io_Pctrl_isPackbt,
  output         io_Pctrl_isPacktb,
  output         io_Pctrl_isPacktt,
  output         io_Pctrl_isPack,
  output [7:0]   io_Pctrl_isSub,
  output         io_Pctrl_isAdder,
  output         io_Pctrl_SrcSigned,
  output         io_Pctrl_Saturating,
  output         io_Pctrl_Translation,
  output         io_Pctrl_LessEqual,
  output         io_Pctrl_LessThan,
  output [79:0]  io_Pctrl_adderRes_ori,
  output [63:0]  io_Pctrl_adderRes,
  output [79:0]  io_Pctrl_adderRes_ori_drophighestbit,
  output         io_Pctrl_Round,
  output         io_Pctrl_ShiftSigned,
  output         io_Pctrl_Arithmetic,
  output         io_Pctrl_isMul_16,
  output         io_Pctrl_isMul_8,
  output         io_Pctrl_isMSW_3232,
  output         io_Pctrl_isMSW_3216,
  output         io_Pctrl_isS1632,
  output         io_Pctrl_isS1664,
  output         io_Pctrl_is832,
  output         io_Pctrl_is3264,
  output         io_Pctrl_is1664,
  output         io_Pctrl_isQ15orQ31,
  output         io_Pctrl_isC31,
  output         io_Pctrl_isQ15_64ONLY,
  output         io_Pctrl_isQ63_64ONLY,
  output         io_Pctrl_isMul_32_64ONLY,
  output         io_Pctrl_isPMA_64ONLY,
  output [17:0]  io_Pctrl_mulres9_0,
  output [17:0]  io_Pctrl_mulres9_1,
  output [17:0]  io_Pctrl_mulres9_2,
  output [17:0]  io_Pctrl_mulres9_3,
  output [33:0]  io_Pctrl_mulres17_0,
  output [33:0]  io_Pctrl_mulres17_1,
  output [65:0]  io_Pctrl_mulres33_0,
  output [129:0] io_Pctrl_mulres65_0
);
  wire [16:0] MulAdd17_0_io_in_srcs_0; // @[PIDU.scala 292:28]
  wire [16:0] MulAdd17_0_io_in_srcs_1; // @[PIDU.scala 292:28]
  wire [33:0] MulAdd17_0_io_out_result; // @[PIDU.scala 292:28]
  wire [16:0] MulAdd17_1_io_in_srcs_0; // @[PIDU.scala 293:28]
  wire [16:0] MulAdd17_1_io_in_srcs_1; // @[PIDU.scala 293:28]
  wire [33:0] MulAdd17_1_io_out_result; // @[PIDU.scala 293:28]
  wire [32:0] MulAdd33_0_io_in_srcs_0; // @[PIDU.scala 294:28]
  wire [32:0] MulAdd33_0_io_in_srcs_1; // @[PIDU.scala 294:28]
  wire [65:0] MulAdd33_0_io_out_result; // @[PIDU.scala 294:28]
  wire [64:0] MulAdd65_0_io_in_srcs_0; // @[PIDU.scala 295:28]
  wire [64:0] MulAdd65_0_io_in_srcs_1; // @[PIDU.scala 295:28]
  wire [129:0] MulAdd65_0_io_out_result; // @[PIDU.scala 295:28]
  wire [8:0] MulAdd9_0_io_in_srcs_0; // @[PIDU.scala 296:28]
  wire [8:0] MulAdd9_0_io_in_srcs_1; // @[PIDU.scala 296:28]
  wire [17:0] MulAdd9_0_io_out_result; // @[PIDU.scala 296:28]
  wire [8:0] MulAdd9_1_io_in_srcs_0; // @[PIDU.scala 297:28]
  wire [8:0] MulAdd9_1_io_in_srcs_1; // @[PIDU.scala 297:28]
  wire [17:0] MulAdd9_1_io_out_result; // @[PIDU.scala 297:28]
  wire [8:0] MulAdd9_2_io_in_srcs_0; // @[PIDU.scala 298:28]
  wire [8:0] MulAdd9_2_io_in_srcs_1; // @[PIDU.scala 298:28]
  wire [17:0] MulAdd9_2_io_out_result; // @[PIDU.scala 298:28]
  wire [8:0] MulAdd9_3_io_in_srcs_0; // @[PIDU.scala 299:28]
  wire [8:0] MulAdd9_3_io_in_srcs_1; // @[PIDU.scala 299:28]
  wire [17:0] MulAdd9_3_io_out_result; // @[PIDU.scala 299:28]
  wire  _T_1 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h2; // @[PIDU.scala 154:36]
  wire  _T_3 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h0; // @[PIDU.scala 154:61]
  wire  _T_5 = io_DecodeIn_ctrl_funct3 == 3'h1; // @[PIDU.scala 154:84]
  wire  _T_10 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0; // @[PIDU.scala 155:72]
  wire  _T_12 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4; // @[PIDU.scala 155:94]
  wire  _T_13 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4; // @[PIDU.scala 155:80]
  wire  _T_14 = _T_3 & (io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4); // @[PIDU.scala 155:51]
  wire  _T_15 = io_DecodeIn_ctrl_funct3 == 3'h2; // @[PIDU.scala 155:113]
  wire  _T_25 = io_DecodeIn_ctrl_funct3 == 3'h0; // @[PIDU.scala 156:113]
  wire  _T_28 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h4; // @[PIDU.scala 157:43]
  wire  _T_38 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h0; // @[PIDU.scala 158:36]
  wire  _T_40 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h2; // @[PIDU.scala 158:62]
  wire  _T_52 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h1; // @[PIDU.scala 160:36]
  wire  _T_71 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h1; // @[PIDU.scala 164:61]
  wire  _T_82 = _T_71 & _T_13; // @[PIDU.scala 165:51]
  wire  _T_96 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h5; // @[PIDU.scala 167:43]
  wire  _T_108 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h3; // @[PIDU.scala 168:62]
  wire  _T_133 = _T_40 & _T_13; // @[PIDU.scala 172:52]
  wire  _T_143 = _T_108 & _T_13; // @[PIDU.scala 173:52]
  wire  _T_166 = io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16; // @[PIDU.scala 176:41]
  wire  _T_170 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h3; // @[PIDU.scala 178:38]
  wire  _T_172 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h5; // @[PIDU.scala 178:63]
  wire  _T_173 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h3 | io_DecodeIn_ctrl_fuOpType[6:4] == 3'h5; // @[PIDU.scala 178:50]
  wire  _T_213 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h6; // @[PIDU.scala 184:44]
  wire  _T_223 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h7; // @[PIDU.scala 185:44]
  wire  _T_234 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h4; // @[PIDU.scala 188:40]
  wire  _T_236 = io_DecodeIn_ctrl_fuOpType[2:1] == 2'h0; // @[PIDU.scala 188:61]
  wire  _T_243 = io_DecodeIn_ctrl_fuOpType[2:1] == 2'h2; // @[PIDU.scala 189:61]
  wire  _T_255 = io_DecodeIn_cf_instr[6:0] == 7'h33; // @[PIDU.scala 190:130]
  wire  _T_258 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h9; // @[PIDU.scala 191:41]
  wire  _T_275 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h1; // @[PIDU.scala 196:35]
  wire  _T_277 = io_DecodeIn_ctrl_fuOpType[4:3] != 2'h0; // @[PIDU.scala 196:56]
  wire  _T_278 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h1 & io_DecodeIn_ctrl_fuOpType[4:3] != 2'h0; // @[PIDU.scala 196:43]
  wire  _T_295 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5; // @[PIDU.scala 198:35]
  wire  _T_297 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6; // @[PIDU.scala 198:56]
  wire  _T_298 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6; // @[PIDU.scala 198:43]
  wire  _T_301 = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6) & _T_108; // @[PIDU.scala 198:64]
  wire  _T_340 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h8; // @[PIDU.scala 202:81]
  wire  _T_341 = _T_278 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h8; // @[PIDU.scala 202:68]
  wire  _T_371 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h3; // @[PIDU.scala 205:35]
  wire  _T_385 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h2; // @[PIDU.scala 207:38]
  wire  _T_387 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hd; // @[PIDU.scala 207:64]
  wire  _T_390 = io_DecodeIn_ctrl_fuOpType[2:1] == 2'h1; // @[PIDU.scala 207:91]
  wire  _T_399 = io_DecodeIn_ctrl_funct3 == 3'h5; // @[PIDU.scala 209:76]
  wire  _T_431 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h7; // @[PIDU.scala 215:37]
  wire  _T_439 = io_DecodeIn_ctrl_fuOpType == 7'h56; // @[PIDU.scala 218:32]
  wire  _T_466 = io_DecodeIn_ctrl_fuOpType == 7'h57; // @[PIDU.scala 224:32]
  wire  _T_530 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'he & (_T_108 | _T_243) & _T_25; // @[PIDU.scala 235:105]
  wire  _T_556 = io_DecodeIn_ctrl_funct3 == 3'h4; // @[PIDU.scala 242:59]
  wire  _T_624 = io_DecodeIn_ctrl_fuOpType == 7'h27; // @[PIDU.scala 252:168]
  wire  _T_633 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hc; // @[PIDU.scala 254:37]
  wire  _T_635 = io_DecodeIn_ctrl_fuOpType[2:0] != 3'h7; // @[PIDU.scala 254:64]
  wire  _T_711 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h1; // @[PIDU.scala 261:72]
  wire  _T_747 = io_DecodeIn_ctrl_fuOpType[1:0] == 2'h1 | _T_258; // @[PIDU.scala 264:57]
  wire [15:0] _GEN_0 = _T_747 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 279:23 281:29]
  wire [15:0] _GEN_1 = _T_747 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 279:23 283:29]
  wire [15:0] _GEN_2 = _T_747 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 279:23 281:29]
  wire [15:0] _GEN_3 = _T_747 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 279:23 283:29]
  wire [63:0] _T_758 = {_GEN_3,_GEN_2,_GEN_1,_GEN_0}; // @[Cat.scala 30:58]
  wire  _T_760 = io_DecodeIn_ctrl_fuOpType[1:0] == 2'h3; // @[PIDU.scala 265:44]
  wire  _T_762 = io_DecodeIn_ctrl_fuOpType[6:3] != 4'hb; // @[PIDU.scala 263:44]
  wire [16:0] _T_765 = {io_DecodeIn_data_src1[15],io_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _T_766 = {1'h0,io_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_4 = _T_762 ? _T_765 : _T_766; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_771 = {io_DecodeIn_data_src1[31],io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _T_772 = {1'h0,io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_5 = _T_762 ? _T_771 : _T_772; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_778 = io_DecodeIn_data_src1[47] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_779 = {_T_778,io_DecodeIn_data_src1[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _T_780 = {17'h0,io_DecodeIn_data_src1[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_6 = _T_762 ? _T_779 : _T_780; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_786 = io_DecodeIn_data_src1[63] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_787 = {_T_786,io_DecodeIn_data_src1[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _T_788 = {49'h0,io_DecodeIn_data_src1[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_7 = _T_762 ? _T_787 : _T_788; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_793 = {_T_758[15],_T_758[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _T_794 = {1'h0,_T_758[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_8 = _T_762 ? _T_793 : _T_794; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_799 = {_T_758[31],_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _T_800 = {1'h0,_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_9 = _T_762 ? _T_799 : _T_800; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_806 = _T_758[47] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_807 = {_T_806,_T_758[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _T_808 = {17'h0,_T_758[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_10 = _T_762 ? _T_807 : _T_808; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_814 = _T_758[63] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_815 = {_T_814,_T_758[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _T_816 = {49'h0,_T_758[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_11 = _T_762 ? _T_815 : _T_816; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_856 = io_DecodeIn_data_src1[31] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_857 = {_T_856,io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _T_858 = {49'h0,io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_17 = _T_762 ? _T_857 : _T_858; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_870 = _T_758[31] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_871 = {_T_870,_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _T_872 = {49'h0,_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_19 = _T_762 ? _T_871 : _T_872; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _GEN_22 = _T_760 ? _GEN_4 : _GEN_4; // @[PIDU.scala 314:35 315:42 328:42]
  wire [16:0] _GEN_23 = _T_760 ? _GEN_5 : 17'h0; // @[PIDU.scala 302:22 314:35 316:42]
  wire [32:0] _GEN_24 = _T_760 ? _GEN_6 : 33'h0; // @[PIDU.scala 303:22 314:35 317:42]
  wire [64:0] _GEN_25 = _T_760 ? _GEN_7 : _GEN_17; // @[PIDU.scala 314:35 318:42 329:42]
  wire [16:0] _GEN_26 = _T_760 ? _GEN_8 : _GEN_8; // @[PIDU.scala 314:35 319:42 330:42]
  wire [16:0] _GEN_27 = _T_760 ? _GEN_9 : 17'h0; // @[PIDU.scala 302:22 314:35 320:42]
  wire [32:0] _GEN_28 = _T_760 ? _GEN_10 : 33'h0; // @[PIDU.scala 303:22 314:35 321:42]
  wire [64:0] _GEN_29 = _T_760 ? _GEN_11 : _GEN_19; // @[PIDU.scala 314:35 322:42 331:42]
  wire [7:0] _GEN_34 = _T_747 ? io_DecodeIn_data_src2[15:8] : io_DecodeIn_data_src2[7:0]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_35 = _T_747 ? io_DecodeIn_data_src2[7:0] : io_DecodeIn_data_src2[15:8]; // @[PIDU.scala 279:23 283:29]
  wire [7:0] _GEN_36 = _T_747 ? io_DecodeIn_data_src2[31:24] : io_DecodeIn_data_src2[23:16]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_37 = _T_747 ? io_DecodeIn_data_src2[23:16] : io_DecodeIn_data_src2[31:24]; // @[PIDU.scala 279:23 283:29]
  wire [7:0] _GEN_38 = _T_747 ? io_DecodeIn_data_src2[47:40] : io_DecodeIn_data_src2[39:32]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_39 = _T_747 ? io_DecodeIn_data_src2[39:32] : io_DecodeIn_data_src2[47:40]; // @[PIDU.scala 279:23 283:29]
  wire [7:0] _GEN_40 = _T_747 ? io_DecodeIn_data_src2[63:56] : io_DecodeIn_data_src2[55:48]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_41 = _T_747 ? io_DecodeIn_data_src2[55:48] : io_DecodeIn_data_src2[63:56]; // @[PIDU.scala 279:23 283:29]
  wire [63:0] _T_914 = {_GEN_41,_GEN_40,_GEN_39,_GEN_38,_GEN_37,_GEN_36,_GEN_35,_GEN_34}; // @[Cat.scala 30:58]
  wire [8:0] _T_921 = {io_DecodeIn_data_src1[7],io_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _T_922 = {1'h0,io_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_42 = _T_762 ? _T_921 : _T_922; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_927 = {io_DecodeIn_data_src1[15],io_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _T_928 = {1'h0,io_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_43 = _T_762 ? _T_927 : _T_928; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_933 = {io_DecodeIn_data_src1[23],io_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _T_934 = {1'h0,io_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_44 = _T_762 ? _T_933 : _T_934; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_939 = {io_DecodeIn_data_src1[31],io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _T_940 = {1'h0,io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_45 = _T_762 ? _T_939 : _T_940; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_946 = io_DecodeIn_data_src1[39] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_947 = {_T_946,io_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _T_948 = {9'h0,io_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_46 = _T_762 ? _T_947 : _T_948; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_954 = io_DecodeIn_data_src1[47] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_955 = {_T_954,io_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _T_956 = {9'h0,io_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_47 = _T_762 ? _T_955 : _T_956; // @[PIDU.scala 268:24 269:15 271:15]
  wire [24:0] _T_962 = io_DecodeIn_data_src1[55] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_963 = {_T_962,io_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _T_964 = {25'h0,io_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_48 = _T_762 ? _T_963 : _T_964; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_970 = io_DecodeIn_data_src1[63] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_971 = {_T_970,io_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _T_972 = {57'h0,io_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_49 = _T_762 ? _T_971 : _T_972; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_977 = {_T_914[7],_T_914[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _T_978 = {1'h0,_T_914[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_50 = _T_762 ? _T_977 : _T_978; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_983 = {_T_914[15],_T_914[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _T_984 = {1'h0,_T_914[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_51 = _T_762 ? _T_983 : _T_984; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_989 = {_T_914[23],_T_914[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _T_990 = {1'h0,_T_914[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_52 = _T_762 ? _T_989 : _T_990; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_995 = {_T_914[31],_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _T_996 = {1'h0,_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_53 = _T_762 ? _T_995 : _T_996; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1002 = _T_914[39] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1003 = {_T_1002,_T_914[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1004 = {9'h0,_T_914[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_54 = _T_762 ? _T_1003 : _T_1004; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1010 = _T_914[47] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1011 = {_T_1010,_T_914[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1012 = {9'h0,_T_914[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_55 = _T_762 ? _T_1011 : _T_1012; // @[PIDU.scala 268:24 269:15 271:15]
  wire [24:0] _T_1018 = _T_914[55] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1019 = {_T_1018,_T_914[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1020 = {25'h0,_T_914[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_56 = _T_762 ? _T_1019 : _T_1020; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1026 = _T_914[63] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1027 = {_T_1026,_T_914[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1028 = {57'h0,_T_914[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_57 = _T_762 ? _T_1027 : _T_1028; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1108 = io_DecodeIn_data_src1[31] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1109 = {_T_1108,io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1110 = {57'h0,io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_69 = _T_762 ? _T_1109 : _T_1110; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1134 = _T_914[31] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1135 = {_T_1134,_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1136 = {57'h0,_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_73 = _T_762 ? _T_1135 : _T_1136; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_78 = _T_760 ? _GEN_42 : _GEN_42; // @[PIDU.scala 338:35 339:42 364:42]
  wire [8:0] _GEN_79 = _T_760 ? _GEN_43 : _GEN_43; // @[PIDU.scala 338:35 340:42 365:42]
  wire [8:0] _GEN_80 = _T_760 ? _GEN_44 : _GEN_44; // @[PIDU.scala 338:35 341:42 366:42]
  wire [8:0] _GEN_81 = _T_760 ? _GEN_45 : 9'h0; // @[PIDU.scala 308:22 338:35 342:42]
  wire [16:0] _GEN_82 = _T_760 ? _GEN_46 : 17'h0; // @[PIDU.scala 301:22 338:35 343:42]
  wire [16:0] _GEN_83 = _T_760 ? _GEN_47 : 17'h0; // @[PIDU.scala 302:22 338:35 344:42]
  wire [32:0] _GEN_84 = _T_760 ? _GEN_48 : 33'h0; // @[PIDU.scala 303:22 338:35 345:42]
  wire [64:0] _GEN_85 = _T_760 ? _GEN_49 : _GEN_69; // @[PIDU.scala 338:35 346:42 367:42]
  wire [8:0] _GEN_86 = _T_760 ? _GEN_50 : _GEN_50; // @[PIDU.scala 338:35 347:42 368:42]
  wire [8:0] _GEN_87 = _T_760 ? _GEN_51 : _GEN_51; // @[PIDU.scala 338:35 348:42 369:42]
  wire [8:0] _GEN_88 = _T_760 ? _GEN_52 : _GEN_52; // @[PIDU.scala 338:35 349:42 370:42]
  wire [8:0] _GEN_89 = _T_760 ? _GEN_53 : 9'h0; // @[PIDU.scala 308:22 338:35 350:42]
  wire [16:0] _GEN_90 = _T_760 ? _GEN_54 : 17'h0; // @[PIDU.scala 301:22 338:35 351:42]
  wire [16:0] _GEN_91 = _T_760 ? _GEN_55 : 17'h0; // @[PIDU.scala 302:22 338:35 352:42]
  wire [32:0] _GEN_92 = _T_760 ? _GEN_56 : 33'h0; // @[PIDU.scala 303:22 338:35 353:42]
  wire [64:0] _GEN_93 = _T_760 ? _GEN_57 : _GEN_73; // @[PIDU.scala 338:35 354:42 371:42]
  wire [32:0] _T_1172 = {io_DecodeIn_data_src1[31],io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1175 = {io_DecodeIn_data_src2[31],io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1181 = io_DecodeIn_data_src1[63] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1182 = {_T_1181,io_DecodeIn_data_src1[63:32]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1186 = io_DecodeIn_data_src2[63] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1187 = {_T_1186,io_DecodeIn_data_src2[63:32]}; // @[Cat.scala 30:58]
  wire  _T_1197 = _T_371 | _T_172 | _T_431; // @[PIDU.scala 388:81]
  wire [15:0] _T_1203 = _T_1197 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 390:52]
  wire [16:0] _T_1206 = _T_1203[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1207 = {_T_1206,_T_1203}; // @[Cat.scala 30:58]
  wire [15:0] _T_1217 = _T_1197 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 393:52]
  wire [48:0] _T_1220 = _T_1217[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1221 = {_T_1220,_T_1217}; // @[Cat.scala 30:58]
  wire  _T_1234 = io_DecodeIn_ctrl_fuOpType[6:3] < 4'h3 | _T_96 & _T_275 & _T_277; // @[PIDU.scala 396:44]
  wire  _T_1239 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h0 | _T_295; // @[PIDU.scala 398:50]
  wire  _T_1244 = _T_711 | _T_297; // @[PIDU.scala 399:50]
  wire [15:0] _T_1248 = _T_1244 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 400:55]
  wire [15:0] _T_1249 = _T_1239 ? io_DecodeIn_data_src1[15:0] : _T_1248; // @[PIDU.scala 400:37]
  wire [15:0] _T_1253 = _T_1244 ? io_DecodeIn_data_src1[47:32] : io_DecodeIn_data_src1[63:48]; // @[PIDU.scala 401:56]
  wire [15:0] _T_1254 = _T_1239 ? io_DecodeIn_data_src1[47:32] : _T_1253; // @[PIDU.scala 401:37]
  wire [15:0] _T_1257 = _T_1239 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 402:37]
  wire [15:0] _T_1260 = _T_1239 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 403:37]
  wire [16:0] _T_1263 = _T_1249[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1264 = {_T_1263,_T_1249}; // @[Cat.scala 30:58]
  wire [16:0] _T_1267 = _T_1257[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1268 = {_T_1267,_T_1257}; // @[Cat.scala 30:58]
  wire [48:0] _T_1273 = _T_1254[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1274 = {_T_1273,_T_1254}; // @[Cat.scala 30:58]
  wire [48:0] _T_1277 = _T_1260[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1278 = {_T_1277,_T_1260}; // @[Cat.scala 30:58]
  wire  _T_1288 = io_DecodeIn_ctrl_fuOpType == 7'h3e; // @[PIDU.scala 411:134]
  wire  _T_1289 = io_DecodeIn_ctrl_fuOpType == 7'h1d | io_DecodeIn_ctrl_fuOpType == 7'h25 | _T_624 |
    io_DecodeIn_ctrl_fuOpType == 7'h3c | io_DecodeIn_ctrl_fuOpType == 7'h3e; // @[PIDU.scala 411:126]
  wire [15:0] _T_1296 = _T_1289 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 413:71]
  wire [15:0] _T_1299 = _T_1289 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 413:105]
  wire [15:0] _T_1302 = _T_1289 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 413:139]
  wire [15:0] _T_1305 = _T_1289 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 413:174]
  wire [16:0] _T_1309 = {_T_1296[15],_T_1296}; // @[Cat.scala 30:58]
  wire [48:0] _T_1318 = _T_1299[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1319 = {_T_1318,_T_1299}; // @[Cat.scala 30:58]
  wire [16:0] _T_1328 = _T_1302[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1329 = {_T_1328,_T_1302}; // @[Cat.scala 30:58]
  wire [48:0] _T_1338 = _T_1305[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1339 = {_T_1338,_T_1305}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_102 = _T_1234 ? _T_1264 : _T_779; // @[PIDU.scala 397:27 404:42 420:42]
  wire [32:0] _GEN_103 = _T_1234 ? _T_1268 : _T_1329; // @[PIDU.scala 397:27 405:42 421:42]
  wire [64:0] _GEN_105 = _T_1234 ? _T_1274 : _T_787; // @[PIDU.scala 397:27 407:42 423:42]
  wire [64:0] _GEN_106 = _T_1234 ? _T_1278 : _T_1339; // @[PIDU.scala 397:27 408:42 424:42]
  wire [16:0] _GEN_108 = _T_1234 ? 17'h0 : _T_765; // @[PIDU.scala 301:22 397:27 414:42]
  wire [16:0] _GEN_109 = _T_1234 ? 17'h0 : _T_1309; // @[PIDU.scala 301:22 397:27 415:42]
  wire [64:0] _GEN_111 = _T_1234 ? 65'h0 : _T_857; // @[PIDU.scala 302:22 397:27 417:42]
  wire [64:0] _GEN_112 = _T_1234 ? 65'h0 : _T_1319; // @[PIDU.scala 302:22 397:27 418:42]
  wire [16:0] _T_1345 = io_DecodeIn_data_src2[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1346 = {_T_1345,io_DecodeIn_data_src2[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1350 = io_DecodeIn_data_src2[31] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1351 = {_T_1350,io_DecodeIn_data_src2[31:16]}; // @[Cat.scala 30:58]
  wire [48:0] _T_1357 = io_DecodeIn_data_src2[47] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1358 = {_T_1357,io_DecodeIn_data_src2[47:32]}; // @[Cat.scala 30:58]
  wire [48:0] _T_1362 = io_DecodeIn_data_src2[63] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1363 = {_T_1362,io_DecodeIn_data_src2[63:48]}; // @[Cat.scala 30:58]
  wire  _T_1370 = ~_T_213; // @[PIDU.scala 438:50]
  wire [8:0] _GEN_114 = _T_1370 ? _T_921 : _T_922; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_115 = _T_1370 ? _T_927 : _T_928; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_116 = _T_1370 ? _T_933 : _T_934; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_117 = _T_1370 ? _T_939 : _T_940; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _GEN_118 = _T_1370 ? _T_947 : _T_948; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _GEN_119 = _T_1370 ? _T_955 : _T_956; // @[PIDU.scala 268:24 269:15 271:15]
  wire [32:0] _GEN_120 = _T_1370 ? _T_963 : _T_964; // @[PIDU.scala 268:24 269:15 271:15]
  wire [64:0] _GEN_121 = _T_1370 ? _T_971 : _T_972; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1420 = {io_DecodeIn_data_src2[7],io_DecodeIn_data_src2[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1421 = {1'h0,io_DecodeIn_data_src2[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_122 = _T_28 ? _T_1420 : _T_1421; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1424 = {io_DecodeIn_data_src2[15],io_DecodeIn_data_src2[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1425 = {1'h0,io_DecodeIn_data_src2[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_123 = _T_28 ? _T_1424 : _T_1425; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1428 = {io_DecodeIn_data_src2[23],io_DecodeIn_data_src2[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1429 = {1'h0,io_DecodeIn_data_src2[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_124 = _T_28 ? _T_1428 : _T_1429; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1432 = {io_DecodeIn_data_src2[31],io_DecodeIn_data_src2[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1433 = {1'h0,io_DecodeIn_data_src2[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_125 = _T_28 ? _T_1432 : _T_1433; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1437 = io_DecodeIn_data_src2[39] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1438 = {_T_1437,io_DecodeIn_data_src2[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1439 = {9'h0,io_DecodeIn_data_src2[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_126 = _T_28 ? _T_1438 : _T_1439; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1443 = io_DecodeIn_data_src2[47] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1444 = {_T_1443,io_DecodeIn_data_src2[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1445 = {9'h0,io_DecodeIn_data_src2[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_127 = _T_28 ? _T_1444 : _T_1445; // @[PIDU.scala 268:24 269:15 271:15]
  wire [24:0] _T_1449 = io_DecodeIn_data_src2[55] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1450 = {_T_1449,io_DecodeIn_data_src2[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1451 = {25'h0,io_DecodeIn_data_src2[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_128 = _T_28 ? _T_1450 : _T_1451; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1455 = io_DecodeIn_data_src2[63] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1456 = {_T_1455,io_DecodeIn_data_src2[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1457 = {57'h0,io_DecodeIn_data_src2[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_129 = _T_28 ? _T_1456 : _T_1457; // @[PIDU.scala 268:24 269:15 271:15]
  wire  _T_1460 = ~io_DecodeIn_ctrl_fuOpType[4]; // @[PIDU.scala 464:30]
  wire [32:0] _T_1464 = {1'h0,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_130 = _T_1460 ? _T_1172 : _T_1464; // @[PIDU.scala 268:24 269:15 271:15]
  wire [64:0] _T_1470 = {33'h0,io_DecodeIn_data_src1[63:32]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_131 = _T_1460 ? _T_1182 : _T_1470; // @[PIDU.scala 268:24 269:15 271:15]
  wire [32:0] _T_1474 = {1'h0,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_132 = _T_1460 ? _T_1175 : _T_1474; // @[PIDU.scala 268:24 269:15 271:15]
  wire [64:0] _T_1480 = {33'h0,io_DecodeIn_data_src2[63:32]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_133 = _T_1460 ? _T_1187 : _T_1480; // @[PIDU.scala 268:24 269:15 271:15]
  wire  _T_1484 = io_DecodeIn_ctrl_fuOpType[4:3] == 2'h0; // @[PIDU.scala 474:36]
  wire  _T_1486 = io_DecodeIn_ctrl_fuOpType[4:3] == 2'h1; // @[PIDU.scala 475:36]
  wire [15:0] _T_1490 = _T_1486 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 476:55]
  wire [15:0] _T_1491 = _T_1484 ? io_DecodeIn_data_src1[15:0] : _T_1490; // @[PIDU.scala 476:37]
  wire [15:0] _T_1495 = _T_1486 ? io_DecodeIn_data_src1[47:32] : io_DecodeIn_data_src1[63:48]; // @[PIDU.scala 477:56]
  wire [15:0] _T_1496 = _T_1484 ? io_DecodeIn_data_src1[47:32] : _T_1495; // @[PIDU.scala 477:37]
  wire [15:0] _T_1499 = _T_1484 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 478:37]
  wire [15:0] _T_1502 = _T_1484 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 479:37]
  wire [16:0] _T_1505 = _T_1491[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1506 = {_T_1505,_T_1491}; // @[Cat.scala 30:58]
  wire [16:0] _T_1509 = _T_1499[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1510 = {_T_1509,_T_1499}; // @[Cat.scala 30:58]
  wire [48:0] _T_1515 = _T_1496[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1516 = {_T_1515,_T_1496}; // @[Cat.scala 30:58]
  wire [48:0] _T_1519 = _T_1502[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1520 = {_T_1519,_T_1502}; // @[Cat.scala 30:58]
  wire  _T_1527 = io_DecodeIn_ctrl_fuOpType == 7'h55 | io_DecodeIn_ctrl_fuOpType == 7'h4e | io_DecodeIn_ctrl_fuOpType
     == 7'h5e; // @[PIDU.scala 487:76]
  wire [15:0] _T_1534 = _T_1527 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 489:71]
  wire [15:0] _T_1537 = _T_1527 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 489:105]
  wire [15:0] _T_1540 = _T_1527 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 489:139]
  wire [15:0] _T_1543 = _T_1527 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 489:174]
  wire [16:0] _T_1547 = {_T_1534[15],_T_1534}; // @[Cat.scala 30:58]
  wire [48:0] _T_1556 = _T_1537[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1557 = {_T_1556,_T_1537}; // @[Cat.scala 30:58]
  wire [16:0] _T_1566 = _T_1540[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1567 = {_T_1566,_T_1540}; // @[Cat.scala 30:58]
  wire [48:0] _T_1576 = _T_1543[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1577 = {_T_1576,_T_1543}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_134 = _T_28 ? _T_1506 : _T_779; // @[PIDU.scala 473:27 480:42 496:42]
  wire [32:0] _GEN_135 = _T_28 ? _T_1510 : _T_1567; // @[PIDU.scala 473:27 481:42 497:42]
  wire [64:0] _GEN_137 = _T_28 ? _T_1516 : _T_787; // @[PIDU.scala 473:27 483:42 499:42]
  wire [64:0] _GEN_138 = _T_28 ? _T_1520 : _T_1577; // @[PIDU.scala 473:27 484:42 500:42]
  wire [16:0] _GEN_140 = _T_28 ? 17'h0 : _T_765; // @[PIDU.scala 301:22 473:27 490:42]
  wire [16:0] _GEN_141 = _T_28 ? 17'h0 : _T_1547; // @[PIDU.scala 301:22 473:27 491:42]
  wire [64:0] _GEN_143 = _T_28 ? 65'h0 : _T_857; // @[PIDU.scala 302:22 473:27 493:42]
  wire [64:0] _GEN_144 = _T_28 ? 65'h0 : _T_1557; // @[PIDU.scala 302:22 473:27 494:42]
  wire  _T_1586 = _T_71 ? _T_1486 : _T_1484; // @[PIDU.scala 505:25]
  wire  _T_1588 = io_DecodeIn_ctrl_fuOpType[4:3] == 2'h2; // @[PIDU.scala 506:48]
  wire  _T_1591 = _T_71 ? io_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 : _T_1486; // @[PIDU.scala 506:25]
  wire [15:0] _T_1595 = _T_1591 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 507:51]
  wire [15:0] _T_1596 = _T_1586 ? io_DecodeIn_data_src1[15:0] : _T_1595; // @[PIDU.scala 507:33]
  wire [15:0] _T_1599 = _T_1586 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 508:33]
  wire [48:0] _T_1602 = _T_1596[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1603 = {_T_1602,_T_1596}; // @[Cat.scala 30:58]
  wire [48:0] _T_1606 = _T_1599[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1607 = {_T_1606,_T_1599}; // @[Cat.scala 30:58]
  wire  _T_1611 = io_DecodeIn_ctrl_fuOpType[6:3] != 4'hf; // @[PIDU.scala 513:59]
  wire [32:0] _T_1615 = io_DecodeIn_data_src1[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1616 = {_T_1615,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1617 = {33'h0,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_146 = _T_1611 ? _T_1616 : _T_1617; // @[PIDU.scala 268:24 269:15 271:15]
  wire [32:0] _T_1623 = io_DecodeIn_data_src2[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1624 = {_T_1623,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1625 = {33'h0,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_147 = _T_1611 ? _T_1624 : _T_1625; // @[PIDU.scala 268:24 269:15 271:15]
  wire [15:0] _T_1635 = _T_1588 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 519:51]
  wire [15:0] _T_1636 = _T_1486 ? io_DecodeIn_data_src1[15:0] : _T_1635; // @[PIDU.scala 519:33]
  wire [15:0] _T_1640 = _T_1588 ? io_DecodeIn_data_src1[47:32] : io_DecodeIn_data_src1[63:48]; // @[PIDU.scala 520:52]
  wire [15:0] _T_1641 = _T_1486 ? io_DecodeIn_data_src1[47:32] : _T_1640; // @[PIDU.scala 520:33]
  wire [15:0] _T_1644 = _T_1486 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 521:33]
  wire [15:0] _T_1647 = _T_1486 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 522:33]
  wire [16:0] _T_1650 = _T_1636[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1651 = {_T_1650,_T_1636}; // @[Cat.scala 30:58]
  wire [16:0] _T_1654 = _T_1644[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1655 = {_T_1654,_T_1644}; // @[Cat.scala 30:58]
  wire [48:0] _T_1660 = _T_1641[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1661 = {_T_1660,_T_1641}; // @[Cat.scala 30:58]
  wire [48:0] _T_1664 = _T_1647[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1665 = {_T_1664,_T_1647}; // @[Cat.scala 30:58]
  wire [31:0] _T_1672 = _T_1486 ? io_DecodeIn_data_src1[31:0] : io_DecodeIn_data_src1[63:32]; // @[PIDU.scala 531:32]
  wire [32:0] _T_1676 = _T_1672[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1677 = {_T_1676,_T_1672}; // @[Cat.scala 30:58]
  wire [31:0] _T_1691 = _T_1588 ? io_DecodeIn_data_src1[31:0] : io_DecodeIn_data_src1[63:32]; // @[PIDU.scala 539:50]
  wire [31:0] _T_1692 = _T_1486 ? io_DecodeIn_data_src1[31:0] : _T_1691; // @[PIDU.scala 539:32]
  wire [31:0] _T_1695 = _T_1486 ? io_DecodeIn_data_src2[31:0] : io_DecodeIn_data_src2[63:32]; // @[PIDU.scala 540:32]
  wire [32:0] _T_1698 = _T_1692[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1699 = {_T_1698,_T_1692}; // @[Cat.scala 30:58]
  wire [32:0] _T_1702 = _T_1695[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1703 = {_T_1702,_T_1695}; // @[Cat.scala 30:58]
  wire  _T_1712 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h7; // @[PIDU.scala 545:87]
  wire  _T_1713 = _T_96 | _T_223 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h7; // @[PIDU.scala 545:74]
  wire [31:0] _T_1718 = _T_1713 ? io_DecodeIn_data_src2[63:32] : io_DecodeIn_data_src2[31:0]; // @[PIDU.scala 548:33]
  wire [31:0] _T_1721 = _T_1713 ? io_DecodeIn_data_src2[31:0] : io_DecodeIn_data_src2[63:32]; // @[PIDU.scala 549:33]
  wire [32:0] _T_1725 = {_T_1718[31],_T_1718}; // @[Cat.scala 30:58]
  wire [32:0] _T_1734 = _T_1721[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1735 = {_T_1734,_T_1721}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_148 = io_Pctrl_isPMA_64ONLY ? _T_1172 : 33'h0; // @[PIDU.scala 303:22 544:42 550:38]
  wire [32:0] _GEN_149 = io_Pctrl_isPMA_64ONLY ? _T_1725 : 33'h0; // @[PIDU.scala 303:22 544:42 551:38]
  wire [64:0] _GEN_151 = io_Pctrl_isPMA_64ONLY ? _T_1182 : 65'h0; // @[PIDU.scala 304:22 544:42 553:38]
  wire [64:0] _GEN_152 = io_Pctrl_isPMA_64ONLY ? _T_1735 : 65'h0; // @[PIDU.scala 304:22 544:42 554:38]
  wire [64:0] _GEN_154 = io_Pctrl_isQ63_64ONLY ? _T_1699 : _GEN_151; // @[PIDU.scala 536:42 541:38]
  wire [64:0] _GEN_155 = io_Pctrl_isQ63_64ONLY ? _T_1703 : _GEN_152; // @[PIDU.scala 536:42 542:38]
  wire [32:0] _GEN_157 = io_Pctrl_isQ63_64ONLY ? 33'h0 : _GEN_148; // @[PIDU.scala 303:22 536:42]
  wire [32:0] _GEN_158 = io_Pctrl_isQ63_64ONLY ? 33'h0 : _GEN_149; // @[PIDU.scala 303:22 536:42]
  wire [64:0] _GEN_160 = io_Pctrl_isMul_32_64ONLY ? _T_1677 : _GEN_154; // @[PIDU.scala 529:45 533:38]
  wire [64:0] _GEN_161 = io_Pctrl_isMul_32_64ONLY ? _T_1187 : _GEN_155; // @[PIDU.scala 529:45 534:38]
  wire [32:0] _GEN_163 = io_Pctrl_isMul_32_64ONLY ? 33'h0 : _GEN_157; // @[PIDU.scala 303:22 529:45]
  wire [32:0] _GEN_164 = io_Pctrl_isMul_32_64ONLY ? 33'h0 : _GEN_158; // @[PIDU.scala 303:22 529:45]
  wire [32:0] _GEN_166 = io_Pctrl_isQ15_64ONLY ? _T_1651 : _GEN_163; // @[PIDU.scala 516:42 523:38]
  wire [32:0] _GEN_167 = io_Pctrl_isQ15_64ONLY ? _T_1655 : _GEN_164; // @[PIDU.scala 516:42 524:38]
  wire [64:0] _GEN_169 = io_Pctrl_isQ15_64ONLY ? _T_1661 : _GEN_160; // @[PIDU.scala 516:42 526:38]
  wire [64:0] _GEN_170 = io_Pctrl_isQ15_64ONLY ? _T_1665 : _GEN_161; // @[PIDU.scala 516:42 527:38]
  wire [64:0] _GEN_172 = io_Pctrl_isC31 ? _GEN_146 : _GEN_169; // @[PIDU.scala 512:35 513:38]
  wire [64:0] _GEN_173 = io_Pctrl_isC31 ? _GEN_147 : _GEN_170; // @[PIDU.scala 512:35 514:38]
  wire [32:0] _GEN_175 = io_Pctrl_isC31 ? 33'h0 : _GEN_166; // @[PIDU.scala 303:22 512:35]
  wire [32:0] _GEN_176 = io_Pctrl_isC31 ? 33'h0 : _GEN_167; // @[PIDU.scala 303:22 512:35]
  wire [64:0] _GEN_178 = io_Pctrl_isQ15orQ31 ? _T_1603 : _GEN_172; // @[PIDU.scala 503:40 509:38]
  wire [64:0] _GEN_179 = io_Pctrl_isQ15orQ31 ? _T_1607 : _GEN_173; // @[PIDU.scala 503:40 510:38]
  wire [32:0] _GEN_181 = io_Pctrl_isQ15orQ31 ? 33'h0 : _GEN_175; // @[PIDU.scala 303:22 503:40]
  wire [32:0] _GEN_182 = io_Pctrl_isQ15orQ31 ? 33'h0 : _GEN_176; // @[PIDU.scala 303:22 503:40]
  wire [32:0] _GEN_184 = io_Pctrl_is1664 ? _GEN_134 : _GEN_181; // @[PIDU.scala 471:36]
  wire [32:0] _GEN_185 = io_Pctrl_is1664 ? _GEN_135 : _GEN_182; // @[PIDU.scala 471:36]
  wire [64:0] _GEN_187 = io_Pctrl_is1664 ? _GEN_137 : _GEN_178; // @[PIDU.scala 471:36]
  wire [64:0] _GEN_188 = io_Pctrl_is1664 ? _GEN_138 : _GEN_179; // @[PIDU.scala 471:36]
  wire [16:0] _GEN_190 = io_Pctrl_is1664 ? _GEN_140 : 17'h0; // @[PIDU.scala 301:22 471:36]
  wire [16:0] _GEN_191 = io_Pctrl_is1664 ? _GEN_141 : 17'h0; // @[PIDU.scala 301:22 471:36]
  wire [64:0] _GEN_193 = io_Pctrl_is1664 ? _GEN_143 : 65'h0; // @[PIDU.scala 302:22 471:36]
  wire [64:0] _GEN_194 = io_Pctrl_is1664 ? _GEN_144 : 65'h0; // @[PIDU.scala 302:22 471:36]
  wire [32:0] _GEN_196 = io_Pctrl_is3264 ? _GEN_130 : _GEN_184; // @[PIDU.scala 462:36 465:38]
  wire [64:0] _GEN_197 = io_Pctrl_is3264 ? _GEN_131 : _GEN_187; // @[PIDU.scala 462:36 466:38]
  wire [32:0] _GEN_198 = io_Pctrl_is3264 ? _GEN_132 : _GEN_185; // @[PIDU.scala 462:36 467:38]
  wire [64:0] _GEN_199 = io_Pctrl_is3264 ? _GEN_133 : _GEN_188; // @[PIDU.scala 462:36 468:38]
  wire [16:0] _GEN_202 = io_Pctrl_is3264 ? 17'h0 : _GEN_190; // @[PIDU.scala 301:22 462:36]
  wire [16:0] _GEN_203 = io_Pctrl_is3264 ? 17'h0 : _GEN_191; // @[PIDU.scala 301:22 462:36]
  wire [64:0] _GEN_205 = io_Pctrl_is3264 ? 65'h0 : _GEN_193; // @[PIDU.scala 302:22 462:36]
  wire [64:0] _GEN_206 = io_Pctrl_is3264 ? 65'h0 : _GEN_194; // @[PIDU.scala 302:22 462:36]
  wire [8:0] _GEN_208 = io_Pctrl_is832 ? _GEN_114 : 9'h0; // @[PIDU.scala 305:22 434:35 438:38]
  wire [8:0] _GEN_209 = io_Pctrl_is832 ? _GEN_115 : 9'h0; // @[PIDU.scala 306:22 434:35 439:38]
  wire [8:0] _GEN_210 = io_Pctrl_is832 ? _GEN_116 : 9'h0; // @[PIDU.scala 307:22 434:35 440:38]
  wire [8:0] _GEN_211 = io_Pctrl_is832 ? _GEN_117 : 9'h0; // @[PIDU.scala 308:22 434:35 441:38]
  wire [16:0] _GEN_212 = io_Pctrl_is832 ? _GEN_118 : _GEN_202; // @[PIDU.scala 434:35 442:38]
  wire [64:0] _GEN_213 = io_Pctrl_is832 ? {{48'd0}, _GEN_119} : _GEN_205; // @[PIDU.scala 434:35 443:38]
  wire [32:0] _GEN_214 = io_Pctrl_is832 ? _GEN_120 : _GEN_196; // @[PIDU.scala 434:35 444:38]
  wire [64:0] _GEN_215 = io_Pctrl_is832 ? _GEN_121 : _GEN_197; // @[PIDU.scala 434:35 445:38]
  wire [8:0] _GEN_216 = io_Pctrl_is832 ? _GEN_122 : 9'h0; // @[PIDU.scala 305:22 434:35 446:38]
  wire [8:0] _GEN_217 = io_Pctrl_is832 ? _GEN_123 : 9'h0; // @[PIDU.scala 306:22 434:35 447:38]
  wire [8:0] _GEN_218 = io_Pctrl_is832 ? _GEN_124 : 9'h0; // @[PIDU.scala 307:22 434:35 448:38]
  wire [8:0] _GEN_219 = io_Pctrl_is832 ? _GEN_125 : 9'h0; // @[PIDU.scala 308:22 434:35 449:38]
  wire [16:0] _GEN_220 = io_Pctrl_is832 ? _GEN_126 : _GEN_203; // @[PIDU.scala 434:35 450:38]
  wire [64:0] _GEN_221 = io_Pctrl_is832 ? {{48'd0}, _GEN_127} : _GEN_206; // @[PIDU.scala 434:35 451:38]
  wire [32:0] _GEN_222 = io_Pctrl_is832 ? _GEN_128 : _GEN_198; // @[PIDU.scala 434:35 452:38]
  wire [64:0] _GEN_223 = io_Pctrl_is832 ? _GEN_129 : _GEN_199; // @[PIDU.scala 434:35 453:38]
  wire [32:0] _GEN_232 = io_Pctrl_isS1664 ? _T_1346 : _GEN_214; // @[PIDU.scala 427:37 428:38]
  wire [32:0] _GEN_233 = io_Pctrl_isS1664 ? _T_1351 : _GEN_222; // @[PIDU.scala 427:37 429:38]
  wire [64:0] _GEN_235 = io_Pctrl_isS1664 ? _T_1358 : _GEN_215; // @[PIDU.scala 427:37 431:38]
  wire [64:0] _GEN_236 = io_Pctrl_isS1664 ? _T_1363 : _GEN_223; // @[PIDU.scala 427:37 432:38]
  wire [8:0] _GEN_238 = io_Pctrl_isS1664 ? 9'h0 : _GEN_208; // @[PIDU.scala 305:22 427:37]
  wire [8:0] _GEN_239 = io_Pctrl_isS1664 ? 9'h0 : _GEN_209; // @[PIDU.scala 306:22 427:37]
  wire [8:0] _GEN_240 = io_Pctrl_isS1664 ? 9'h0 : _GEN_210; // @[PIDU.scala 307:22 427:37]
  wire [8:0] _GEN_241 = io_Pctrl_isS1664 ? 9'h0 : _GEN_211; // @[PIDU.scala 308:22 427:37]
  wire [16:0] _GEN_242 = io_Pctrl_isS1664 ? 17'h0 : _GEN_212; // @[PIDU.scala 301:22 427:37]
  wire [64:0] _GEN_243 = io_Pctrl_isS1664 ? 65'h0 : _GEN_213; // @[PIDU.scala 302:22 427:37]
  wire [8:0] _GEN_244 = io_Pctrl_isS1664 ? 9'h0 : _GEN_216; // @[PIDU.scala 305:22 427:37]
  wire [8:0] _GEN_245 = io_Pctrl_isS1664 ? 9'h0 : _GEN_217; // @[PIDU.scala 306:22 427:37]
  wire [8:0] _GEN_246 = io_Pctrl_isS1664 ? 9'h0 : _GEN_218; // @[PIDU.scala 307:22 427:37]
  wire [8:0] _GEN_247 = io_Pctrl_isS1664 ? 9'h0 : _GEN_219; // @[PIDU.scala 308:22 427:37]
  wire [16:0] _GEN_248 = io_Pctrl_isS1664 ? 17'h0 : _GEN_220; // @[PIDU.scala 301:22 427:37]
  wire [64:0] _GEN_249 = io_Pctrl_isS1664 ? 65'h0 : _GEN_221; // @[PIDU.scala 302:22 427:37]
  wire [32:0] _GEN_256 = io_Pctrl_isS1632 ? _GEN_102 : _GEN_232; // @[PIDU.scala 395:37]
  wire [32:0] _GEN_257 = io_Pctrl_isS1632 ? _GEN_103 : _GEN_233; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_259 = io_Pctrl_isS1632 ? _GEN_105 : _GEN_235; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_260 = io_Pctrl_isS1632 ? _GEN_106 : _GEN_236; // @[PIDU.scala 395:37]
  wire [16:0] _GEN_262 = io_Pctrl_isS1632 ? _GEN_108 : _GEN_242; // @[PIDU.scala 395:37]
  wire [16:0] _GEN_263 = io_Pctrl_isS1632 ? _GEN_109 : _GEN_248; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_265 = io_Pctrl_isS1632 ? _GEN_111 : _GEN_243; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_266 = io_Pctrl_isS1632 ? _GEN_112 : _GEN_249; // @[PIDU.scala 395:37]
  wire [8:0] _GEN_268 = io_Pctrl_isS1632 ? 9'h0 : _GEN_238; // @[PIDU.scala 305:22 395:37]
  wire [8:0] _GEN_269 = io_Pctrl_isS1632 ? 9'h0 : _GEN_239; // @[PIDU.scala 306:22 395:37]
  wire [8:0] _GEN_270 = io_Pctrl_isS1632 ? 9'h0 : _GEN_240; // @[PIDU.scala 307:22 395:37]
  wire [8:0] _GEN_271 = io_Pctrl_isS1632 ? 9'h0 : _GEN_241; // @[PIDU.scala 308:22 395:37]
  wire [8:0] _GEN_272 = io_Pctrl_isS1632 ? 9'h0 : _GEN_244; // @[PIDU.scala 305:22 395:37]
  wire [8:0] _GEN_273 = io_Pctrl_isS1632 ? 9'h0 : _GEN_245; // @[PIDU.scala 306:22 395:37]
  wire [8:0] _GEN_274 = io_Pctrl_isS1632 ? 9'h0 : _GEN_246; // @[PIDU.scala 307:22 395:37]
  wire [8:0] _GEN_275 = io_Pctrl_isS1632 ? 9'h0 : _GEN_247; // @[PIDU.scala 308:22 395:37]
  wire [32:0] _GEN_280 = io_Pctrl_isMSW_3216 ? _T_1172 : _GEN_256; // @[PIDU.scala 386:40 389:38]
  wire [32:0] _GEN_281 = io_Pctrl_isMSW_3216 ? _T_1207 : _GEN_257; // @[PIDU.scala 386:40 390:38]
  wire [64:0] _GEN_283 = io_Pctrl_isMSW_3216 ? _T_1182 : _GEN_259; // @[PIDU.scala 386:40 392:38]
  wire [64:0] _GEN_284 = io_Pctrl_isMSW_3216 ? _T_1221 : _GEN_260; // @[PIDU.scala 386:40 393:38]
  wire [16:0] _GEN_286 = io_Pctrl_isMSW_3216 ? 17'h0 : _GEN_262; // @[PIDU.scala 301:22 386:40]
  wire [16:0] _GEN_287 = io_Pctrl_isMSW_3216 ? 17'h0 : _GEN_263; // @[PIDU.scala 301:22 386:40]
  wire [64:0] _GEN_289 = io_Pctrl_isMSW_3216 ? 65'h0 : _GEN_265; // @[PIDU.scala 302:22 386:40]
  wire [64:0] _GEN_290 = io_Pctrl_isMSW_3216 ? 65'h0 : _GEN_266; // @[PIDU.scala 302:22 386:40]
  wire [8:0] _GEN_292 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_268; // @[PIDU.scala 305:22 386:40]
  wire [8:0] _GEN_293 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_269; // @[PIDU.scala 306:22 386:40]
  wire [8:0] _GEN_294 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_270; // @[PIDU.scala 307:22 386:40]
  wire [8:0] _GEN_295 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_271; // @[PIDU.scala 308:22 386:40]
  wire [8:0] _GEN_296 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_272; // @[PIDU.scala 305:22 386:40]
  wire [8:0] _GEN_297 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_273; // @[PIDU.scala 306:22 386:40]
  wire [8:0] _GEN_298 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_274; // @[PIDU.scala 307:22 386:40]
  wire [8:0] _GEN_299 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_275; // @[PIDU.scala 308:22 386:40]
  wire [32:0] _GEN_304 = io_Pctrl_isMSW_3232 ? _T_1172 : _GEN_280; // @[PIDU.scala 378:40 380:38]
  wire [32:0] _GEN_305 = io_Pctrl_isMSW_3232 ? _T_1175 : _GEN_281; // @[PIDU.scala 378:40 381:38]
  wire [64:0] _GEN_307 = io_Pctrl_isMSW_3232 ? _T_1182 : _GEN_283; // @[PIDU.scala 378:40 383:38]
  wire [64:0] _GEN_308 = io_Pctrl_isMSW_3232 ? _T_1187 : _GEN_284; // @[PIDU.scala 378:40 384:38]
  wire [16:0] _GEN_310 = io_Pctrl_isMSW_3232 ? 17'h0 : _GEN_286; // @[PIDU.scala 301:22 378:40]
  wire [16:0] _GEN_311 = io_Pctrl_isMSW_3232 ? 17'h0 : _GEN_287; // @[PIDU.scala 301:22 378:40]
  wire [64:0] _GEN_313 = io_Pctrl_isMSW_3232 ? 65'h0 : _GEN_289; // @[PIDU.scala 302:22 378:40]
  wire [64:0] _GEN_314 = io_Pctrl_isMSW_3232 ? 65'h0 : _GEN_290; // @[PIDU.scala 302:22 378:40]
  wire [8:0] _GEN_316 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_292; // @[PIDU.scala 305:22 378:40]
  wire [8:0] _GEN_317 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_293; // @[PIDU.scala 306:22 378:40]
  wire [8:0] _GEN_318 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_294; // @[PIDU.scala 307:22 378:40]
  wire [8:0] _GEN_319 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_295; // @[PIDU.scala 308:22 378:40]
  wire [8:0] _GEN_320 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_296; // @[PIDU.scala 305:22 378:40]
  wire [8:0] _GEN_321 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_297; // @[PIDU.scala 306:22 378:40]
  wire [8:0] _GEN_322 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_298; // @[PIDU.scala 307:22 378:40]
  wire [8:0] _GEN_323 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_299; // @[PIDU.scala 308:22 378:40]
  wire [8:0] _GEN_328 = io_Pctrl_isMul_8 ? _GEN_78 : _GEN_316; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_329 = io_Pctrl_isMul_8 ? _GEN_79 : _GEN_317; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_330 = io_Pctrl_isMul_8 ? _GEN_80 : _GEN_318; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_331 = io_Pctrl_isMul_8 ? _GEN_81 : _GEN_319; // @[PIDU.scala 335:37]
  wire [16:0] _GEN_332 = io_Pctrl_isMul_8 ? _GEN_82 : _GEN_310; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_333 = io_Pctrl_isMul_8 ? {{48'd0}, _GEN_83} : _GEN_313; // @[PIDU.scala 335:37]
  wire [32:0] _GEN_334 = io_Pctrl_isMul_8 ? _GEN_84 : _GEN_304; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_335 = io_Pctrl_isMul_8 ? _GEN_85 : _GEN_307; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_336 = io_Pctrl_isMul_8 ? _GEN_86 : _GEN_320; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_337 = io_Pctrl_isMul_8 ? _GEN_87 : _GEN_321; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_338 = io_Pctrl_isMul_8 ? _GEN_88 : _GEN_322; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_339 = io_Pctrl_isMul_8 ? _GEN_89 : _GEN_323; // @[PIDU.scala 335:37]
  wire [16:0] _GEN_340 = io_Pctrl_isMul_8 ? _GEN_90 : _GEN_311; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_341 = io_Pctrl_isMul_8 ? {{48'd0}, _GEN_91} : _GEN_314; // @[PIDU.scala 335:37]
  wire [32:0] _GEN_342 = io_Pctrl_isMul_8 ? _GEN_92 : _GEN_305; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_343 = io_Pctrl_isMul_8 ? _GEN_93 : _GEN_308; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_353 = io_Pctrl_isMul_16 ? {{48'd0}, _GEN_23} : _GEN_333; // @[PIDU.scala 311:32]
  wire [64:0] _GEN_357 = io_Pctrl_isMul_16 ? {{48'd0}, _GEN_27} : _GEN_341; // @[PIDU.scala 311:32]
  wire  _T_1748 = io_Pctrl_isSub_64 | io_Pctrl_isSub_32 | io_Pctrl_isSub_16 | io_Pctrl_isSub_8 | io_Pctrl_isComp_16; // @[PIDU.scala 633:87]
  wire [1:0] _GEN_376 = io_Pctrl_isCrsa_32 | io_Pctrl_isStsa_32 ? 2'h2 : 2'h0; // @[PIDU.scala 632:20 642:56 643:23]
  wire [1:0] _GEN_377 = io_Pctrl_isCras_32 | io_Pctrl_isStas_32 ? 2'h1 : _GEN_376; // @[PIDU.scala 640:56 641:23]
  wire [3:0] _GEN_378 = io_Pctrl_isCrsa_16 | io_Pctrl_isStsa_16 ? 4'ha : {{2'd0}, _GEN_377}; // @[PIDU.scala 638:56 639:23]
  wire [3:0] _GEN_379 = io_Pctrl_isCras_16 | io_Pctrl_isStas_16 ? 4'h5 : _GEN_378; // @[PIDU.scala 636:56 637:23]
  wire  _T_1775 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hb; // @[PIDU.scala 648:104]
  wire  _T_1781 = ~io_Pctrl_isSt; // @[PIDU.scala 649:29]
  wire  _T_1787 = ~io_DecodeIn_ctrl_fuOpType[3]; // @[PIDU.scala 649:82]
  wire  _T_1804 = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8; // @[PIDU.scala 797:32]
  wire  _T_1811 = io_Pctrl_isPbs ? 1'h0 : io_Pctrl_SrcSigned; // @[PIDU.scala 798:74]
  wire  _T_1812 = io_Pctrl_isMaxMin_8 ? _T_1787 : _T_1811; // @[PIDU.scala 798:34]
  wire [8:0] _T_1817 = {{1'd0}, io_DecodeIn_data_src1[7:0]}; // @[PIDU.scala 671:57]
  wire  _GEN_384 = _T_1812 & _T_1817[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1831 = {{1'd0}, io_DecodeIn_data_src1[15:8]}; // @[PIDU.scala 671:57]
  wire  _GEN_388 = _T_1812 & _T_1831[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1845 = {{1'd0}, io_DecodeIn_data_src1[23:16]}; // @[PIDU.scala 671:57]
  wire  _GEN_392 = _T_1812 & _T_1845[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1859 = {{1'd0}, io_DecodeIn_data_src1[31:24]}; // @[PIDU.scala 671:57]
  wire  _GEN_396 = _T_1812 & _T_1859[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1873 = {{1'd0}, io_DecodeIn_data_src1[39:32]}; // @[PIDU.scala 671:57]
  wire  _GEN_400 = _T_1812 & _T_1873[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1887 = {{1'd0}, io_DecodeIn_data_src1[47:40]}; // @[PIDU.scala 671:57]
  wire  _GEN_404 = _T_1812 & _T_1887[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1901 = {{1'd0}, io_DecodeIn_data_src1[55:48]}; // @[PIDU.scala 671:57]
  wire  _GEN_408 = _T_1812 & _T_1901[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1915 = {{1'd0}, io_DecodeIn_data_src1[63:56]}; // @[PIDU.scala 671:57]
  wire  _GEN_412 = _T_1812 & _T_1915[7]; // @[PIDU.scala 673:28]
  wire [30:0] _T_1933 = {1'h0,_GEN_412,_T_1915[7:0],1'h0,_GEN_408,_T_1901[7:0],1'h0,_GEN_404,_T_1887[7:0],1'h0}; // @[Cat.scala 30:58]
  wire [60:0] _T_1942 = {_T_1933,_GEN_400,_T_1873[7:0],1'h0,_GEN_396,_T_1859[7:0],1'h0,_GEN_392,_T_1845[7:0],1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_1947 = {_T_1942,_GEN_388,_T_1831[7:0],1'h0,_GEN_384,_T_1817[7:0]}; // @[Cat.scala 30:58]
  wire [7:0] _T_1952 = io_Pctrl_isSub[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1953 = io_DecodeIn_data_src2[7:0] ^ _T_1952; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_577 = {{7'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_1956 = _T_1953 + _GEN_577; // @[PIDU.scala 671:57]
  wire  _T_1962 = io_Pctrl_isSub[0] & _T_1956 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_414 = io_Pctrl_isSub[0] & _T_1956 == 8'h80 ? 1'h0 : _T_1956[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_1965 = io_Pctrl_isSub[0] & _T_1956 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_416 = _T_1812 ? _GEN_414 : _T_1965; // @[PIDU.scala 673:28]
  wire [7:0] _T_1971 = io_Pctrl_isSub[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1972 = io_DecodeIn_data_src2[15:8] ^ _T_1971; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_578 = {{7'd0}, io_Pctrl_isSub[1]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_1975 = _T_1972 + _GEN_578; // @[PIDU.scala 671:57]
  wire  _T_1981 = io_Pctrl_isSub[1] & _T_1975 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_418 = io_Pctrl_isSub[1] & _T_1975 == 8'h80 ? 1'h0 : _T_1975[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_1984 = io_Pctrl_isSub[1] & _T_1975 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_420 = _T_1812 ? _GEN_418 : _T_1984; // @[PIDU.scala 673:28]
  wire [7:0] _T_1990 = io_Pctrl_isSub[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1991 = io_DecodeIn_data_src2[23:16] ^ _T_1990; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_579 = {{7'd0}, io_Pctrl_isSub[2]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_1994 = _T_1991 + _GEN_579; // @[PIDU.scala 671:57]
  wire  _T_2000 = io_Pctrl_isSub[2] & _T_1994 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_422 = io_Pctrl_isSub[2] & _T_1994 == 8'h80 ? 1'h0 : _T_1994[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2003 = io_Pctrl_isSub[2] & _T_1994 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_424 = _T_1812 ? _GEN_422 : _T_2003; // @[PIDU.scala 673:28]
  wire [7:0] _T_2009 = io_Pctrl_isSub[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2010 = io_DecodeIn_data_src2[31:24] ^ _T_2009; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_580 = {{7'd0}, io_Pctrl_isSub[3]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2013 = _T_2010 + _GEN_580; // @[PIDU.scala 671:57]
  wire  _T_2019 = io_Pctrl_isSub[3] & _T_2013 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_426 = io_Pctrl_isSub[3] & _T_2013 == 8'h80 ? 1'h0 : _T_2013[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2022 = io_Pctrl_isSub[3] & _T_2013 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_428 = _T_1812 ? _GEN_426 : _T_2022; // @[PIDU.scala 673:28]
  wire [7:0] _T_2028 = io_Pctrl_isSub[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2029 = io_DecodeIn_data_src2[39:32] ^ _T_2028; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_581 = {{7'd0}, io_Pctrl_isSub[4]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2032 = _T_2029 + _GEN_581; // @[PIDU.scala 671:57]
  wire  _T_2038 = io_Pctrl_isSub[4] & _T_2032 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_430 = io_Pctrl_isSub[4] & _T_2032 == 8'h80 ? 1'h0 : _T_2032[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2041 = io_Pctrl_isSub[4] & _T_2032 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_432 = _T_1812 ? _GEN_430 : _T_2041; // @[PIDU.scala 673:28]
  wire [7:0] _T_2047 = io_Pctrl_isSub[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2048 = io_DecodeIn_data_src2[47:40] ^ _T_2047; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_582 = {{7'd0}, io_Pctrl_isSub[5]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2051 = _T_2048 + _GEN_582; // @[PIDU.scala 671:57]
  wire  _T_2057 = io_Pctrl_isSub[5] & _T_2051 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_434 = io_Pctrl_isSub[5] & _T_2051 == 8'h80 ? 1'h0 : _T_2051[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2060 = io_Pctrl_isSub[5] & _T_2051 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_436 = _T_1812 ? _GEN_434 : _T_2060; // @[PIDU.scala 673:28]
  wire [7:0] _T_2066 = io_Pctrl_isSub[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2067 = io_DecodeIn_data_src2[55:48] ^ _T_2066; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_583 = {{7'd0}, io_Pctrl_isSub[6]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2070 = _T_2067 + _GEN_583; // @[PIDU.scala 671:57]
  wire  _T_2076 = io_Pctrl_isSub[6] & _T_2070 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_438 = io_Pctrl_isSub[6] & _T_2070 == 8'h80 ? 1'h0 : _T_2070[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2079 = io_Pctrl_isSub[6] & _T_2070 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_440 = _T_1812 ? _GEN_438 : _T_2079; // @[PIDU.scala 673:28]
  wire [7:0] _T_2085 = io_Pctrl_isSub[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2086 = io_DecodeIn_data_src2[63:56] ^ _T_2085; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_584 = {{7'd0}, io_Pctrl_isSub[7]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2089 = _T_2086 + _GEN_584; // @[PIDU.scala 671:57]
  wire  _T_2095 = io_Pctrl_isSub[7] & _T_2089 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_442 = io_Pctrl_isSub[7] & _T_2089 == 8'h80 ? 1'h0 : _T_2089[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2098 = io_Pctrl_isSub[7] & _T_2089 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_444 = _T_1812 ? _GEN_442 : _T_2098; // @[PIDU.scala 673:28]
  wire [30:0] _T_2108 = {1'h0,_GEN_444,_T_2089,1'h0,_GEN_440,_T_2070,1'h0,_GEN_436,_T_2051,1'h0}; // @[Cat.scala 30:58]
  wire [60:0] _T_2117 = {_T_2108,_GEN_432,_T_2032,1'h0,_GEN_428,_T_2013,1'h0,_GEN_424,_T_1994,1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_2122 = {_T_2117,_GEN_420,_T_1975,1'h0,_GEN_416,_T_1956}; // @[Cat.scala 30:58]
  wire [29:0] _T_2221 = {3'h0,_T_1915[6:0],1'h0,1'h0,1'h0,_T_1901[6:0],1'h0,1'h0,1'h0,_T_1887[6:0]}; // @[Cat.scala 30:58]
  wire [50:0] _T_2230 = {_T_2221,1'h0,1'h0,1'h0,_T_1873[6:0],1'h0,1'h0,1'h0,_T_1859[6:0],1'h0}; // @[Cat.scala 30:58]
  wire [71:0] _T_2239 = {_T_2230,1'h0,1'h0,_T_1845[6:0],1'h0,1'h0,1'h0,_T_1831[6:0],1'h0,1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_2241 = {_T_2239,1'h0,_T_1817[6:0]}; // @[Cat.scala 30:58]
  wire [22:0] _T_2371 = {2'h0,_T_2095,_T_2089[6:0],1'h0,1'h0,_T_2076,_T_2070[6:0],1'h0,1'h0,_T_2057}; // @[Cat.scala 30:58]
  wire [49:0] _T_2380 = {_T_2371,_T_2051[6:0],1'h0,1'h0,_T_2038,_T_2032[6:0],1'h0,1'h0,_T_2019,_T_2013[6:0]}; // @[Cat.scala 30:58]
  wire [70:0] _T_2389 = {_T_2380,1'h0,1'h0,_T_2000,_T_1994[6:0],1'h0,1'h0,_T_1981,_T_1975[6:0],1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_2392 = {_T_2389,1'h0,_T_1962,_T_1956[6:0]}; // @[Cat.scala 30:58]
  wire  _T_2395 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16; // @[PIDU.scala 803:81]
  wire  _T_2402 = io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15; // @[PIDU.scala 804:51]
  wire [63:0] _T_2405 = {48'h0,io_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2406 = io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15 ? _T_2405 : io_DecodeIn_data_src1; // @[PIDU.scala 804:31]
  wire [63:0] _T_2410 = {48'h0,io_DecodeIn_data_src2[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2411 = _T_2402 ? _T_2410 : io_DecodeIn_data_src2; // @[PIDU.scala 805:31]
  wire  _T_2417 = io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15 ? _T_1787 : io_Pctrl_SrcSigned; // @[PIDU.scala 806:34]
  wire [16:0] _T_2424 = {{1'd0}, _T_2406[15:0]}; // @[PIDU.scala 671:57]
  wire  _GEN_480 = _T_2417 & _T_2424[15]; // @[PIDU.scala 673:28]
  wire [16:0] _T_2438 = {{1'd0}, _T_2406[31:16]}; // @[PIDU.scala 671:57]
  wire  _GEN_484 = _T_2417 & _T_2438[15]; // @[PIDU.scala 673:28]
  wire [16:0] _T_2452 = {{1'd0}, _T_2406[47:32]}; // @[PIDU.scala 671:57]
  wire  _GEN_488 = _T_2417 & _T_2452[15]; // @[PIDU.scala 673:28]
  wire [16:0] _T_2466 = {{1'd0}, _T_2406[63:48]}; // @[PIDU.scala 671:57]
  wire  _GEN_492 = _T_2417 & _T_2466[15]; // @[PIDU.scala 673:28]
  wire [54:0] _T_2484 = {1'h0,_GEN_492,_T_2466[15:0],1'h0,_GEN_488,_T_2452[15:0],1'h0,_GEN_484,_T_2438[15:0],1'h0}; // @[Cat.scala 30:58]
  wire [71:0] _T_2486 = {_T_2484,_GEN_480,_T_2424[15:0]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_493 = _T_166 ? _T_2411[31:16] : _T_2411[15:0]; // @[PIDU.scala 663:21 664:23 666:29]
  wire [15:0] _T_2491 = io_Pctrl_isSub[0] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2492 = _GEN_493 ^ _T_2491; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_593 = {{15'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2495 = _T_2492 + _GEN_593; // @[PIDU.scala 671:57]
  wire  _T_2501 = io_Pctrl_isSub[0] & _T_2495 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_494 = io_Pctrl_isSub[0] & _T_2495 == 16'h8000 ? 1'h0 : _T_2495[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2504 = io_Pctrl_isSub[0] & _T_2495 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_496 = _T_2417 ? _GEN_494 : _T_2504; // @[PIDU.scala 673:28]
  wire [15:0] _GEN_497 = _T_166 ? _T_2411[15:0] : _T_2411[31:16]; // @[PIDU.scala 663:21 664:23 668:29]
  wire [15:0] _T_2510 = io_Pctrl_isSub[1] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2511 = _GEN_497 ^ _T_2510; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_594 = {{15'd0}, io_Pctrl_isSub[1]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2514 = _T_2511 + _GEN_594; // @[PIDU.scala 671:57]
  wire  _T_2520 = io_Pctrl_isSub[1] & _T_2514 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_498 = io_Pctrl_isSub[1] & _T_2514 == 16'h8000 ? 1'h0 : _T_2514[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2523 = io_Pctrl_isSub[1] & _T_2514 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_500 = _T_2417 ? _GEN_498 : _T_2523; // @[PIDU.scala 673:28]
  wire [15:0] _GEN_501 = _T_166 ? _T_2411[63:48] : _T_2411[47:32]; // @[PIDU.scala 663:21 664:23 666:29]
  wire [15:0] _T_2529 = io_Pctrl_isSub[2] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2530 = _GEN_501 ^ _T_2529; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_595 = {{15'd0}, io_Pctrl_isSub[2]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2533 = _T_2530 + _GEN_595; // @[PIDU.scala 671:57]
  wire  _T_2539 = io_Pctrl_isSub[2] & _T_2533 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_502 = io_Pctrl_isSub[2] & _T_2533 == 16'h8000 ? 1'h0 : _T_2533[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2542 = io_Pctrl_isSub[2] & _T_2533 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_504 = _T_2417 ? _GEN_502 : _T_2542; // @[PIDU.scala 673:28]
  wire [15:0] _GEN_505 = _T_166 ? _T_2411[47:32] : _T_2411[63:48]; // @[PIDU.scala 663:21 664:23 668:29]
  wire [15:0] _T_2548 = io_Pctrl_isSub[3] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2549 = _GEN_505 ^ _T_2548; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_596 = {{15'd0}, io_Pctrl_isSub[3]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2552 = _T_2549 + _GEN_596; // @[PIDU.scala 671:57]
  wire  _T_2558 = io_Pctrl_isSub[3] & _T_2552 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_506 = io_Pctrl_isSub[3] & _T_2552 == 16'h8000 ? 1'h0 : _T_2552[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2561 = io_Pctrl_isSub[3] & _T_2552 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_508 = _T_2417 ? _GEN_506 : _T_2561; // @[PIDU.scala 673:28]
  wire [54:0] _T_2571 = {1'h0,_GEN_508,_T_2552,1'h0,_GEN_504,_T_2533,1'h0,_GEN_500,_T_2514,1'h0}; // @[Cat.scala 30:58]
  wire [71:0] _T_2573 = {_T_2571,_GEN_496,_T_2495}; // @[Cat.scala 30:58]
  wire [53:0] _T_2628 = {3'h0,_T_2466[14:0],1'h0,1'h0,1'h0,_T_2452[14:0],1'h0,1'h0,1'h0,_T_2438[14:0]}; // @[Cat.scala 30:58]
  wire [71:0] _T_2632 = {_T_2628,1'h0,1'h0,1'h0,_T_2424[14:0]}; // @[Cat.scala 30:58]
  wire [38:0] _T_2702 = {2'h0,_T_2558,_T_2552[14:0],1'h0,1'h0,_T_2539,_T_2533[14:0],1'h0,1'h0,_T_2520}; // @[Cat.scala 30:58]
  wire [71:0] _T_2707 = {_T_2702,_T_2514[14:0],1'h0,1'h0,_T_2501,_T_2495[14:0]}; // @[Cat.scala 30:58]
  wire  _T_2710 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32; // @[PIDU.scala 812:81]
  wire  _T_2720 = io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31; // @[PIDU.scala 813:93]
  wire [63:0] _T_2723 = {32'h0,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2724 = io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2723 :
    io_DecodeIn_data_src1; // @[PIDU.scala 813:31]
  wire [63:0] _T_2730 = {32'h0,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2731 = _T_2720 ? _T_2730 : io_DecodeIn_data_src2; // @[PIDU.scala 814:31]
  wire  _T_2740 = io_Pctrl_isMaxMin_32 ? io_DecodeIn_ctrl_fuOpType[3] : io_Pctrl_SrcSigned; // @[PIDU.scala 815:135]
  wire  _T_2741 = _T_2720 ? _T_1787 : _T_2740; // @[PIDU.scala 815:34]
  wire  _T_2742 = io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32; // @[PIDU.scala 816:50]
  wire [32:0] _T_2748 = {{1'd0}, _T_2724[31:0]}; // @[PIDU.scala 671:57]
  wire  _GEN_528 = _T_2741 & _T_2748[31]; // @[PIDU.scala 673:28]
  wire [32:0] _T_2762 = {{1'd0}, _T_2724[63:32]}; // @[PIDU.scala 671:57]
  wire  _GEN_532 = _T_2741 & _T_2762[31]; // @[PIDU.scala 673:28]
  wire [67:0] _T_2776 = {1'h0,_GEN_532,_T_2762[31:0],1'h0,_GEN_528,_T_2748[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_533 = _T_2742 ? _T_2731[63:32] : _T_2731[31:0]; // @[PIDU.scala 663:21 664:23 666:29]
  wire [31:0] _T_2781 = io_Pctrl_isSub[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2782 = _GEN_533 ^ _T_2781; // @[PIDU.scala 671:32]
  wire [31:0] _GEN_601 = {{31'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [31:0] _T_2785 = _T_2782 + _GEN_601; // @[PIDU.scala 671:57]
  wire  _T_2791 = io_Pctrl_isSub[0] & _T_2785 == 32'h80000000; // @[PIDU.scala 675:31]
  wire  _GEN_534 = io_Pctrl_isSub[0] & _T_2785 == 32'h80000000 ? 1'h0 : _T_2785[31]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2794 = io_Pctrl_isSub[0] & _T_2785 != 32'h0; // @[PIDU.scala 678:31]
  wire  _GEN_536 = _T_2741 ? _GEN_534 : _T_2794; // @[PIDU.scala 673:28]
  wire [31:0] _GEN_537 = _T_2742 ? _T_2731[31:0] : _T_2731[63:32]; // @[PIDU.scala 663:21 664:23 668:29]
  wire [31:0] _T_2800 = io_Pctrl_isSub[1] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2801 = _GEN_537 ^ _T_2800; // @[PIDU.scala 671:32]
  wire [31:0] _GEN_602 = {{31'd0}, io_Pctrl_isSub[1]}; // @[PIDU.scala 671:57]
  wire [31:0] _T_2804 = _T_2801 + _GEN_602; // @[PIDU.scala 671:57]
  wire  _T_2810 = io_Pctrl_isSub[1] & _T_2804 == 32'h80000000; // @[PIDU.scala 675:31]
  wire  _GEN_538 = io_Pctrl_isSub[1] & _T_2804 == 32'h80000000 ? 1'h0 : _T_2804[31]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2813 = io_Pctrl_isSub[1] & _T_2804 != 32'h0; // @[PIDU.scala 678:31]
  wire  _GEN_540 = _T_2741 ? _GEN_538 : _T_2813; // @[PIDU.scala 673:28]
  wire [67:0] _T_2819 = {1'h0,_GEN_540,_T_2804,1'h0,_GEN_536,_T_2785}; // @[Cat.scala 30:58]
  wire [67:0] _T_2848 = {3'h0,_T_2762[30:0],1'h0,1'h0,1'h0,_T_2748[30:0]}; // @[Cat.scala 30:58]
  wire [67:0] _T_2885 = {2'h0,_T_2810,_T_2804[30:0],1'h0,1'h0,_T_2791,_T_2785[30:0]}; // @[Cat.scala 30:58]
  wire  _T_2889 = io_Pctrl_isMaxMin_XLEN | io_Pctrl_isAve | io_Pctrl_SrcSigned; // @[PIDU.scala 822:34]
  wire [64:0] _T_2893 = {{1'd0}, io_DecodeIn_data_src1}; // @[PIDU.scala 671:57]
  wire  _GEN_551 = _T_2889 & _T_2893[63]; // @[PIDU.scala 673:28]
  wire [65:0] _T_2904 = {1'h0,_GEN_551,_T_2893[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2908 = io_Pctrl_isSub[0] ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2909 = io_DecodeIn_data_src2 ^ _T_2908; // @[PIDU.scala 671:32]
  wire [63:0] _GEN_605 = {{63'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [63:0] _T_2912 = _T_2909 + _GEN_605; // @[PIDU.scala 671:57]
  wire  _T_2918 = io_Pctrl_isSub[0] & _T_2912 == 64'h8000000000000000; // @[PIDU.scala 675:31]
  wire  _GEN_552 = io_Pctrl_isSub[0] & _T_2912 == 64'h8000000000000000 ? 1'h0 : _T_2912[63]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2921 = io_Pctrl_isSub[0] & _T_2912 != 64'h0; // @[PIDU.scala 678:31]
  wire  _GEN_554 = _T_2889 ? _GEN_552 : _T_2921; // @[PIDU.scala 673:28]
  wire [65:0] _T_2924 = {1'h0,_GEN_554,_T_2912}; // @[Cat.scala 30:58]
  wire [65:0] _T_2937 = {3'h0,_T_2893[62:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_2954 = {2'h0,_T_2918,_T_2912[62:0]}; // @[Cat.scala 30:58]
  wire [67:0] _GEN_561 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2776 : {{2'd0}, _T_2904}; // @[PIDU.scala 812:251 817:18]
  wire [67:0] _GEN_562 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2819 : {{2'd0}, _T_2924}; // @[PIDU.scala 812:251 818:18]
  wire [67:0] _GEN_563 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2848 : {{2'd0}, _T_2937}; // @[PIDU.scala 812:251 819:33]
  wire [67:0] _GEN_564 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2885 : {{2'd0}, _T_2954}; // @[PIDU.scala 812:251 820:33]
  wire [71:0] _GEN_565 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2486 : {{4'd0}, _GEN_561}; // @[PIDU.scala 803:231 808:18]
  wire [71:0] _GEN_566 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2573 : {{4'd0}, _GEN_562}; // @[PIDU.scala 803:231 809:18]
  wire [71:0] _GEN_567 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2632 : {{4'd0}, _GEN_563}; // @[PIDU.scala 803:231 810:33]
  wire [71:0] _GEN_568 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2707 : {{4'd0}, _GEN_564}; // @[PIDU.scala 803:231 811:33]
  wire [79:0] add1 = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 | io_Pctrl_isPbs ?
    _T_1947 : {{8'd0}, _GEN_565}; // @[PIDU.scala 797:111 799:18]
  wire [79:0] add2 = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 | io_Pctrl_isPbs ?
    _T_2122 : {{8'd0}, _GEN_566}; // @[PIDU.scala 797:111 800:18]
  wire [79:0] add1_drophighestbit = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 |
    io_Pctrl_isPbs ? _T_2241 : {{8'd0}, _GEN_567}; // @[PIDU.scala 797:111 801:33]
  wire [79:0] add2_drophighestbit = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 |
    io_Pctrl_isPbs ? _T_2392 : {{8'd0}, _GEN_568}; // @[PIDU.scala 797:111 802:33]
  wire [80:0] _T_2955 = add1 + add2; // @[PIDU.scala 840:35]
  wire [80:0] _T_2956 = add1_drophighestbit + add2_drophighestbit; // @[PIDU.scala 841:65]
  wire [63:0] _T_2973 = {io_Pctrl_adderRes_ori[77:70],io_Pctrl_adderRes_ori[67:60],io_Pctrl_adderRes_ori[57:50],
    io_Pctrl_adderRes_ori[47:40],io_Pctrl_adderRes_ori[37:30],io_Pctrl_adderRes_ori[27:20],io_Pctrl_adderRes_ori[17:10],
    io_Pctrl_adderRes_ori[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2987 = {io_Pctrl_adderRes_ori[69:54],io_Pctrl_adderRes_ori[51:36],io_Pctrl_adderRes_ori[33:18],
    io_Pctrl_adderRes_ori[15:0]}; // @[Cat.scala 30:58]
  wire  _T_2991 = _T_2710 | io_Pctrl_isAdd_Q31; // @[PIDU.scala 862:98]
  wire [63:0] _T_2999 = {io_Pctrl_adderRes_ori[65:34],io_Pctrl_adderRes_ori[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_574 = _T_2991 | io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 | io_Pctrl_isStas_32 |
    io_Pctrl_isStsa_32 ? _T_2999 : io_Pctrl_adderRes_ori[63:0]; // @[PIDU.scala 863:111 864:27]
  wire [63:0] _GEN_575 = _T_2395 | io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15 | io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 ?
    _T_2987 : _GEN_574; // @[PIDU.scala 860:90 861:27]
  wire  _T_3010 = _T_297 & (~io_DecodeIn_ctrl_fuOpType[1] | _T_760); // @[PIDU.scala 871:54]
  wire  _T_3025 = (_T_3010 | _T_1712 & (_T_236 & io_DecodeIn_ctrl_func24 | _T_243 & io_DecodeIn_ctrl_func23)) & _T_25; // @[PIDU.scala 872:126]
  wire  _T_3030 = _T_297 | _T_340; // @[PIDU.scala 873:63]
  wire  _T_3036 = _T_3025 | (io_Pctrl_isRs_32 & (_T_297 | _T_340) | io_Pctrl_isLR_32 & io_DecodeIn_ctrl_fuOpType[4]); // @[PIDU.scala 873:21]
  wire  _T_3040 = _T_3036 | io_Pctrl_isLR_Q31 & io_DecodeIn_ctrl_fuOpType[3]; // @[PIDU.scala 874:21]
  wire  _T_3041 = _T_3040 | io_Pctrl_isRs_XLEN; // @[PIDU.scala 875:21]
  MulAdd_onestage MulAdd17_0 ( // @[PIDU.scala 292:28]
    .io_in_srcs_0(MulAdd17_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd17_0_io_in_srcs_1),
    .io_out_result(MulAdd17_0_io_out_result)
  );
  MulAdd_onestage MulAdd17_1 ( // @[PIDU.scala 293:28]
    .io_in_srcs_0(MulAdd17_1_io_in_srcs_0),
    .io_in_srcs_1(MulAdd17_1_io_in_srcs_1),
    .io_out_result(MulAdd17_1_io_out_result)
  );
  MulAdd_onestage_2 MulAdd33_0 ( // @[PIDU.scala 294:28]
    .io_in_srcs_0(MulAdd33_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd33_0_io_in_srcs_1),
    .io_out_result(MulAdd33_0_io_out_result)
  );
  MulAdd_onestage_3 MulAdd65_0 ( // @[PIDU.scala 295:28]
    .io_in_srcs_0(MulAdd65_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd65_0_io_in_srcs_1),
    .io_out_result(MulAdd65_0_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_0 ( // @[PIDU.scala 296:28]
    .io_in_srcs_0(MulAdd9_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_0_io_in_srcs_1),
    .io_out_result(MulAdd9_0_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_1 ( // @[PIDU.scala 297:28]
    .io_in_srcs_0(MulAdd9_1_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_1_io_in_srcs_1),
    .io_out_result(MulAdd9_1_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_2 ( // @[PIDU.scala 298:28]
    .io_in_srcs_0(MulAdd9_2_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_2_io_in_srcs_1),
    .io_out_result(MulAdd9_2_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_3 ( // @[PIDU.scala 299:28]
    .io_in_srcs_0(MulAdd9_3_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_3_io_in_srcs_1),
    .io_out_result(MulAdd9_3_io_out_result)
  );
  assign io_Pctrl_isAdd_64 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h2 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h0 &
    io_DecodeIn_ctrl_funct3 == 3'h1; // @[PIDU.scala 154:74]
  assign io_Pctrl_isAdd_32 = _T_3 & (io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4) &
    io_DecodeIn_ctrl_funct3 == 3'h2; // @[PIDU.scala 155:103]
  assign io_Pctrl_isAdd_16 = _T_14 & io_DecodeIn_ctrl_funct3 == 3'h0; // @[PIDU.scala 156:103]
  assign io_Pctrl_isAdd_8 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h4 & _T_13 & _T_25; // @[PIDU.scala 157:103]
  assign io_Pctrl_isAdd_Q15 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h0 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h2 & _T_5; // @[PIDU.scala 158:75]
  assign io_Pctrl_isAdd_Q31 = _T_38 & _T_3 & _T_5; // @[PIDU.scala 159:75]
  assign io_Pctrl_isAdd_C31 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h1 & _T_3 & _T_5; // @[PIDU.scala 160:75]
  assign io_Pctrl_isAve = io_DecodeIn_ctrl_fuOpType == 7'h70 & _T_25; // @[PIDU.scala 161:48]
  assign io_Pctrl_isAdd = io_Pctrl_isAdd_64 | io_Pctrl_isAdd_32 | io_Pctrl_isAdd_16 | io_Pctrl_isAdd_8 |
    io_Pctrl_isAdd_Q15 | io_Pctrl_isAdd_Q31 | io_Pctrl_isAdd_C31 | io_Pctrl_isAve; // @[PIDU.scala 162:163]
  assign io_Pctrl_isSub_64 = _T_1 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h1 & _T_5; // @[PIDU.scala 164:74]
  assign io_Pctrl_isSub_32 = _T_71 & _T_13 & _T_15; // @[PIDU.scala 165:103]
  assign io_Pctrl_isSub_16 = _T_82 & _T_25; // @[PIDU.scala 166:103]
  assign io_Pctrl_isSub_8 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h5 & _T_13 & _T_25; // @[PIDU.scala 167:103]
  assign io_Pctrl_isSub_Q15 = _T_38 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h3 & _T_5; // @[PIDU.scala 168:75]
  assign io_Pctrl_isSub_Q31 = _T_38 & _T_71 & _T_5; // @[PIDU.scala 169:75]
  assign io_Pctrl_isSub_C31 = _T_52 & _T_71 & _T_5; // @[PIDU.scala 170:75]
  assign io_Pctrl_isCras_16 = _T_40 & _T_13 & _T_25; // @[PIDU.scala 172:103]
  assign io_Pctrl_isCrsa_16 = _T_108 & _T_13 & _T_25; // @[PIDU.scala 173:103]
  assign io_Pctrl_isCras_32 = _T_133 & _T_15; // @[PIDU.scala 174:103]
  assign io_Pctrl_isCrsa_32 = _T_143 & _T_15; // @[PIDU.scala 175:103]
  assign io_Pctrl_isCr = io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32; // @[PIDU.scala 176:83]
  assign io_Pctrl_isStas_16 = (io_DecodeIn_ctrl_fuOpType[6:5] == 2'h3 | io_DecodeIn_ctrl_fuOpType[6:4] == 3'h5) & _T_40
     & _T_15; // @[PIDU.scala 178:103]
  assign io_Pctrl_isStsa_16 = _T_173 & _T_108 & _T_15; // @[PIDU.scala 179:103]
  assign io_Pctrl_isStas_32 = _T_173 & _T_3 & _T_15; // @[PIDU.scala 180:103]
  assign io_Pctrl_isStsa_32 = _T_173 & _T_71 & _T_15; // @[PIDU.scala 181:103]
  assign io_Pctrl_isSt = io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isStas_32 | io_Pctrl_isStsa_32; // @[PIDU.scala 182:83]
  assign io_Pctrl_isComp_16 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h6 & _T_13 & _T_25; // @[PIDU.scala 184:96]
  assign io_Pctrl_isComp_8 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h7 & _T_13 & _T_25; // @[PIDU.scala 185:96]
  assign io_Pctrl_isCompare = io_Pctrl_isComp_16 | io_Pctrl_isComp_8; // @[PIDU.scala 186:46]
  assign io_Pctrl_isMaxMin_16 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h4 & io_DecodeIn_ctrl_fuOpType[2:1] == 2'h0 & _T_25; // @[PIDU.scala 188:69]
  assign io_Pctrl_isMaxMin_8 = _T_234 & io_DecodeIn_ctrl_fuOpType[2:1] == 2'h2 & _T_25; // @[PIDU.scala 189:69]
  assign io_Pctrl_isMaxMin_XLEN = io_DecodeIn_ctrl_fuOpType == 7'h5 & io_DecodeIn_ctrl_funct3[2] & ~
    io_DecodeIn_ctrl_funct3[0] & io_DecodeIn_cf_instr[6:0] == 7'h33; // @[PIDU.scala 190:101]
  assign io_Pctrl_isMaxMin_32 = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h9 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'ha) &
    _T_236 & _T_15; // @[PIDU.scala 191:104]
  assign io_Pctrl_isMaxMin = io_Pctrl_isMaxMin_16 | io_Pctrl_isMaxMin_8 | io_Pctrl_isMaxMin_XLEN | io_Pctrl_isMaxMin_32; // @[PIDU.scala 192:98]
  assign io_Pctrl_isPbs = io_DecodeIn_ctrl_fuOpType[6:1] == 6'h3f & _T_25; // @[PIDU.scala 194:53]
  assign io_Pctrl_isRs_16 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h1 & io_DecodeIn_ctrl_fuOpType[4:3] != 2'h0 & _T_236 &
    _T_25; // @[PIDU.scala 196:85]
  assign io_Pctrl_isLs_16 = _T_278 & _T_40 & _T_25; // @[PIDU.scala 197:85]
  assign io_Pctrl_isLR_16 = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6) & _T_108
     & _T_25; // @[PIDU.scala 198:85]
  assign io_Pctrl_isRs_8 = _T_278 & _T_243 & _T_25; // @[PIDU.scala 199:85]
  assign io_Pctrl_isLs_8 = _T_278 & _T_213 & _T_25; // @[PIDU.scala 200:85]
  assign io_Pctrl_isLR_8 = _T_298 & _T_223 & _T_25; // @[PIDU.scala 201:85]
  assign io_Pctrl_isRs_32 = (_T_278 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h8) & _T_236 & _T_15; // @[PIDU.scala 202:111]
  assign io_Pctrl_isLs_32 = _T_341 & _T_40 & _T_15; // @[PIDU.scala 203:111]
  assign io_Pctrl_isLR_32 = _T_301 & _T_15; // @[PIDU.scala 204:86]
  assign io_Pctrl_isLR_Q31 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h3 & _T_223 & _T_5; // @[PIDU.scala 205:74]
  assign io_Pctrl_isLs_Q31 = _T_52 & _T_108 & _T_5; // @[PIDU.scala 206:74]
  assign io_Pctrl_isRs_XLEN = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h2 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'hd) &
    io_DecodeIn_ctrl_fuOpType[2:1] == 2'h1 & _T_5; // @[PIDU.scala 207:103]
  assign io_Pctrl_isSRAIWU = io_DecodeIn_ctrl_fuOpType == 7'h1a & _T_5; // @[PIDU.scala 208:47]
  assign io_Pctrl_isFSRW = io_DecodeIn_cf_instr[26:25] == 2'h2 & io_DecodeIn_ctrl_funct3 == 3'h5 &
    io_DecodeIn_ctrl_fuOpType == 7'h3b; // @[PIDU.scala 209:91]
  assign io_Pctrl_isWext = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h6 & _T_223 & _T_25; // @[PIDU.scala 210:76]
  assign io_Pctrl_isShifter = io_Pctrl_isRs_16 | io_Pctrl_isLs_16 | io_Pctrl_isLR_16 | io_Pctrl_isRs_8 | io_Pctrl_isLs_8
     | io_Pctrl_isLR_8 | io_Pctrl_isRs_32 | io_Pctrl_isLs_32 | io_Pctrl_isLR_32 | io_Pctrl_isLs_Q31 | io_Pctrl_isLR_Q31
     | io_Pctrl_isRs_XLEN | io_Pctrl_isSRAIWU | io_Pctrl_isFSRW | io_Pctrl_isWext; // @[PIDU.scala 211:292]
  assign io_Pctrl_isClip_16 = io_DecodeIn_ctrl_fuOpType == 7'h42 & _T_25; // @[PIDU.scala 213:49]
  assign io_Pctrl_isClip_8 = io_DecodeIn_ctrl_fuOpType == 7'h46 & _T_25; // @[PIDU.scala 214:49]
  assign io_Pctrl_isclip_32 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h7 & _T_40 & _T_25; // @[PIDU.scala 215:75]
  assign io_Pctrl_isClip = io_Pctrl_isClip_16 | io_Pctrl_isClip_8 | io_Pctrl_isclip_32; // @[PIDU.scala 216:66]
  assign io_Pctrl_isSat_16 = io_DecodeIn_ctrl_fuOpType == 7'h56 & io_DecodeIn_data_src2[4:0] == 5'h11 & _T_25; // @[PIDU.scala 218:77]
  assign io_Pctrl_isSat_8 = _T_439 & io_DecodeIn_data_src2[4:0] == 5'h10 & _T_25; // @[PIDU.scala 219:77]
  assign io_Pctrl_isSat_32 = _T_439 & io_DecodeIn_data_src2[4:0] == 5'h12 & _T_25; // @[PIDU.scala 220:77]
  assign io_Pctrl_isSat_W = _T_439 & io_DecodeIn_data_src2[4:0] == 5'h14 & _T_25; // @[PIDU.scala 221:77]
  assign io_Pctrl_isSat = io_Pctrl_isSat_16 | io_Pctrl_isSat_8 | io_Pctrl_isSat_32 | io_Pctrl_isSat_W; // @[PIDU.scala 222:84]
  assign io_Pctrl_isCnt_16 = io_DecodeIn_ctrl_fuOpType == 7'h57 & io_DecodeIn_data_src2[4:1] == 4'h4 & _T_25; // @[PIDU.scala 224:76]
  assign io_Pctrl_isCnt_8 = _T_466 & io_DecodeIn_data_src2[4:1] == 4'h0 & _T_25; // @[PIDU.scala 225:76]
  assign io_Pctrl_isCnt_32 = _T_466 & io_DecodeIn_data_src2[4:1] == 4'hc & _T_25; // @[PIDU.scala 226:76]
  assign io_Pctrl_isCnt = io_Pctrl_isCnt_16 | io_Pctrl_isCnt_8 | io_Pctrl_isCnt_32; // @[PIDU.scala 227:64]
  assign io_Pctrl_isSwap_16 = _T_10 & _T_223 & _T_5; // @[PIDU.scala 229:72]
  assign io_Pctrl_isSwap_8 = _T_439 & (io_DecodeIn_data_src2[4:0] == 5'h18 & _T_25 & io_DecodeIn_cf_instrType == 5'h15
     | io_DecodeIn_data_src2[5:0] == 6'h8 & _T_399 & io_DecodeIn_cf_instrType == 5'h17); // @[PIDU.scala 230:49]
  assign io_Pctrl_isSwap = io_Pctrl_isSwap_16 | io_Pctrl_isSwap_8; // @[PIDU.scala 231:46]
  assign io_Pctrl_isUnpack = _T_439 & (io_DecodeIn_data_src2[4:3] == 2'h1 | io_DecodeIn_data_src2[4:0] == 5'h13 |
    io_DecodeIn_data_src2[4:0] == 5'h17) & _T_25; // @[PIDU.scala 233:132]
  assign io_Pctrl_isBitrev = _T_530 | io_DecodeIn_ctrl_fuOpType == 7'h35 & _T_399 & io_DecodeIn_cf_instr[6:0] == 7'h13
     & io_DecodeIn_data_src2[4:0] == 5'h1f; // @[PIDU.scala 236:24]
  assign io_Pctrl_isCmix = io_DecodeIn_cf_instr[14:12] == 3'h1 & _T_255 & io_DecodeIn_cf_instr[26:25] == 2'h3; // @[PIDU.scala 238:114]
  assign io_Pctrl_isInsertb = _T_439 & io_DecodeIn_cf_instr[24:23] == 2'h0 & _T_25; // @[PIDU.scala 240:92]
  assign io_Pctrl_isPackbb = io_DecodeIn_ctrl_fuOpType == 7'h4 & io_DecodeIn_ctrl_funct3 == 3'h4 & _T_255; // @[PIDU.scala 242:72]
  assign io_Pctrl_isPackbt = io_DecodeIn_ctrl_fuOpType == 7'hf & _T_15; // @[PIDU.scala 243:49]
  assign io_Pctrl_isPacktb = io_DecodeIn_ctrl_fuOpType == 7'h1f & _T_15; // @[PIDU.scala 244:49]
  assign io_Pctrl_isPacktt = io_DecodeIn_ctrl_fuOpType == 7'h24 & _T_556 & _T_255; // @[PIDU.scala 245:72]
  assign io_Pctrl_isPack = io_Pctrl_isPackbb | io_Pctrl_isPackbt | io_Pctrl_isPacktb | io_Pctrl_isPacktt; // @[PIDU.scala 246:85]
  assign io_Pctrl_isSub = _T_1748 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin | io_Pctrl_isPbs | io_Pctrl_isSub_Q15 |
    io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 ? 8'hff : {{4'd0}, _GEN_379}; // @[PIDU.scala 634:125 635:23]
  assign io_Pctrl_isAdder = (io_Pctrl_isSub != 8'h0 | io_Pctrl_isAdd | io_Pctrl_isCr | io_Pctrl_isSt) & ~
    io_Pctrl_isCompare & ~io_Pctrl_isMaxMin & ~io_Pctrl_isPbs; // @[PIDU.scala 646:142]
  assign io_Pctrl_SrcSigned = _T_38 | _T_234 | io_Pctrl_isSt & (io_DecodeIn_ctrl_fuOpType[6:3] == 4'hb | _T_633); // @[PIDU.scala 648:73]
  assign io_Pctrl_Saturating = ~io_Pctrl_isSt & io_DecodeIn_ctrl_fuOpType[3] | io_Pctrl_isSt & ~
    io_DecodeIn_ctrl_fuOpType[3]; // @[PIDU.scala 649:62]
  assign io_Pctrl_Translation = ~io_Pctrl_Saturating & (_T_1781 & ~_T_12 | io_Pctrl_isSt & (_T_1775 | _T_387)); // @[PIDU.scala 650:50]
  assign io_Pctrl_LessEqual = io_Pctrl_Saturating; // @[PIDU.scala 651:26]
  assign io_Pctrl_LessThan = io_Pctrl_Translation; // @[PIDU.scala 652:26]
  assign io_Pctrl_adderRes_ori = _T_2955[79:0]; // @[PIDU.scala 840:27]
  assign io_Pctrl_adderRes = _T_1804 | io_Pctrl_isPbs ? _T_2973 : _GEN_575; // @[PIDU.scala 857:65 858:27]
  assign io_Pctrl_adderRes_ori_drophighestbit = _T_2956[79:0]; // @[PIDU.scala 841:42]
  assign io_Pctrl_Round = _T_3041 | io_Pctrl_isSRAIWU; // @[PIDU.scala 876:21]
  assign io_Pctrl_ShiftSigned = io_Pctrl_isLR_16 | io_Pctrl_isLR_8 | io_Pctrl_isLR_32 | io_Pctrl_isLR_Q31 |
    io_Pctrl_isLs_Q31 | io_Pctrl_isLs_32 & _T_3030 | (io_Pctrl_isLs_16 | io_Pctrl_isLs_8) & (_T_297 |
    io_DecodeIn_ctrl_fuOpType == 7'h3a & io_DecodeIn_ctrl_func24 | _T_1288 & io_DecodeIn_ctrl_func23); // @[PIDU.scala 877:191]
  assign io_Pctrl_Arithmetic = (io_Pctrl_isRs_16 | io_Pctrl_isRs_8 | io_Pctrl_isRs_32) & ~io_DecodeIn_ctrl_fuOpType[0]
     | io_Pctrl_isLR_16 | io_Pctrl_isLR_8 | io_Pctrl_isLR_32 | io_Pctrl_isLR_Q31 | io_Pctrl_isRs_XLEN |
    io_Pctrl_isSRAIWU; // @[PIDU.scala 878:209]
  assign io_Pctrl_isMul_16 = ~io_DecodeIn_ctrl_fuOpType[2] & _T_25; // @[PIDU.scala 248:43]
  assign io_Pctrl_isMul_8 = io_DecodeIn_ctrl_fuOpType[2] & _T_25 & io_DecodeIn_ctrl_fuOpType[6:3] != 4'hc; // @[PIDU.scala 249:61]
  assign io_Pctrl_isMSW_3232 = _T_275 & _T_236 & _T_5; // @[PIDU.scala 250:76]
  assign io_Pctrl_isMSW_3216 = (_T_275 & _T_390 | io_DecodeIn_ctrl_fuOpType[6] & _T_223) & _T_5; // @[PIDU.scala 251:126]
  assign io_Pctrl_isS1632 = ~io_DecodeIn_ctrl_fuOpType[6] & (_T_28 | _T_96 & io_DecodeIn_ctrl_fuOpType[6:3] > 4'h2 |
    _T_213 & io_DecodeIn_ctrl_fuOpType[5] | io_DecodeIn_ctrl_fuOpType == 7'h27) & _T_5; // @[PIDU.scala 252:187]
  assign io_Pctrl_isS1664 = io_DecodeIn_ctrl_fuOpType == 7'h2f & _T_5; // @[PIDU.scala 253:49]
  assign io_Pctrl_is832 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hc & io_DecodeIn_ctrl_fuOpType[2:0] != 3'h7 & _T_25; // @[PIDU.scala 254:77]
  assign io_Pctrl_is3264 = _T_1 & _T_390 & _T_5; // @[PIDU.scala 255:74]
  assign io_Pctrl_is1664 = _T_1 & _T_635 & _T_5; // @[PIDU.scala 256:75]
  assign io_Pctrl_isQ15orQ31 = (_T_10 & (_T_213 | _T_96) | _T_170 & _T_71 & _T_277) & _T_5; // @[PIDU.scala 257:183]
  assign io_Pctrl_isC31 = (_T_431 & _T_3 | _T_633 & _T_390) & _T_5; // @[PIDU.scala 258:130]
  assign io_Pctrl_isQ15_64ONLY = _T_170 & _T_277 & io_DecodeIn_ctrl_fuOpType[2] & io_DecodeIn_ctrl_fuOpType[1:0] != 2'h3
     & _T_5; // @[PIDU.scala 259:123]
  assign io_Pctrl_isQ63_64ONLY = _T_278 & _T_96 & _T_15; // @[PIDU.scala 260:102]
  assign io_Pctrl_isMul_32_64ONLY = (_T_385 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h1) & _T_28 & _T_15; // @[PIDU.scala 261:113]
  assign io_Pctrl_isPMA_64ONLY = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h3 & _T_243 | _T_12 & io_DecodeIn_ctrl_fuOpType[2]
     | (_T_28 | _T_213) & _T_275 & _T_277) & _T_15; // @[PIDU.scala 262:223]
  assign io_Pctrl_mulres9_0 = MulAdd9_0_io_out_result; // @[PIDU.scala 622:25]
  assign io_Pctrl_mulres9_1 = MulAdd9_1_io_out_result; // @[PIDU.scala 623:25]
  assign io_Pctrl_mulres9_2 = MulAdd9_2_io_out_result; // @[PIDU.scala 624:25]
  assign io_Pctrl_mulres9_3 = MulAdd9_3_io_out_result; // @[PIDU.scala 625:25]
  assign io_Pctrl_mulres17_0 = MulAdd17_0_io_out_result; // @[PIDU.scala 626:25]
  assign io_Pctrl_mulres17_1 = MulAdd17_1_io_out_result; // @[PIDU.scala 627:25]
  assign io_Pctrl_mulres33_0 = MulAdd33_0_io_out_result; // @[PIDU.scala 628:25]
  assign io_Pctrl_mulres65_0 = MulAdd65_0_io_out_result; // @[PIDU.scala 629:25]
  assign MulAdd17_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? _GEN_22 : _GEN_332; // @[PIDU.scala 311:32]
  assign MulAdd17_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? _GEN_26 : _GEN_340; // @[PIDU.scala 311:32]
  assign MulAdd17_1_io_in_srcs_0 = _GEN_353[16:0];
  assign MulAdd17_1_io_in_srcs_1 = _GEN_357[16:0];
  assign MulAdd33_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? _GEN_24 : _GEN_334; // @[PIDU.scala 311:32]
  assign MulAdd33_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? _GEN_28 : _GEN_342; // @[PIDU.scala 311:32]
  assign MulAdd65_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? _GEN_25 : _GEN_335; // @[PIDU.scala 311:32]
  assign MulAdd65_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? _GEN_29 : _GEN_343; // @[PIDU.scala 311:32]
  assign MulAdd9_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_328; // @[PIDU.scala 305:22 311:32]
  assign MulAdd9_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_336; // @[PIDU.scala 305:22 311:32]
  assign MulAdd9_1_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_329; // @[PIDU.scala 306:22 311:32]
  assign MulAdd9_1_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_337; // @[PIDU.scala 306:22 311:32]
  assign MulAdd9_2_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_330; // @[PIDU.scala 307:22 311:32]
  assign MulAdd9_2_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_338; // @[PIDU.scala 307:22 311:32]
  assign MulAdd9_3_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_331; // @[PIDU.scala 308:22 311:32]
  assign MulAdd9_3_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_339; // @[PIDU.scala 308:22 311:32]
endmodule
module PIDU_1(
  input  [63:0]  io_DecodeIn_cf_instr,
  input  [4:0]   io_DecodeIn_cf_instrType,
  input  [6:0]   io_DecodeIn_ctrl_fuOpType,
  input  [2:0]   io_DecodeIn_ctrl_funct3,
  input          io_DecodeIn_ctrl_func24,
  input          io_DecodeIn_ctrl_func23,
  input  [63:0]  io_DecodeIn_data_src1,
  input  [63:0]  io_DecodeIn_data_src2,
  output         io_Pctrl_isAdd_64,
  output         io_Pctrl_isAdd_32,
  output         io_Pctrl_isAdd_16,
  output         io_Pctrl_isAdd_8,
  output         io_Pctrl_isAdd_Q15,
  output         io_Pctrl_isAdd_Q31,
  output         io_Pctrl_isAdd_C31,
  output         io_Pctrl_isAve,
  output         io_Pctrl_isAdd,
  output         io_Pctrl_isSub_64,
  output         io_Pctrl_isSub_32,
  output         io_Pctrl_isSub_16,
  output         io_Pctrl_isSub_8,
  output         io_Pctrl_isSub_Q15,
  output         io_Pctrl_isSub_Q31,
  output         io_Pctrl_isSub_C31,
  output         io_Pctrl_isCras_16,
  output         io_Pctrl_isCrsa_16,
  output         io_Pctrl_isCras_32,
  output         io_Pctrl_isCrsa_32,
  output         io_Pctrl_isCr,
  output         io_Pctrl_isStas_16,
  output         io_Pctrl_isStsa_16,
  output         io_Pctrl_isStas_32,
  output         io_Pctrl_isStsa_32,
  output         io_Pctrl_isSt,
  output         io_Pctrl_isComp_16,
  output         io_Pctrl_isComp_8,
  output         io_Pctrl_isCompare,
  output         io_Pctrl_isMaxMin_16,
  output         io_Pctrl_isMaxMin_8,
  output         io_Pctrl_isMaxMin_XLEN,
  output         io_Pctrl_isMaxMin_32,
  output         io_Pctrl_isMaxMin,
  output         io_Pctrl_isPbs,
  output         io_Pctrl_isRs_16,
  output         io_Pctrl_isLs_16,
  output         io_Pctrl_isLR_16,
  output         io_Pctrl_isRs_8,
  output         io_Pctrl_isLs_8,
  output         io_Pctrl_isLR_8,
  output         io_Pctrl_isRs_32,
  output         io_Pctrl_isLs_32,
  output         io_Pctrl_isLR_32,
  output         io_Pctrl_isLR_Q31,
  output         io_Pctrl_isLs_Q31,
  output         io_Pctrl_isRs_XLEN,
  output         io_Pctrl_isSRAIWU,
  output         io_Pctrl_isFSRW,
  output         io_Pctrl_isWext,
  output         io_Pctrl_isShifter,
  output         io_Pctrl_isClip_16,
  output         io_Pctrl_isClip_8,
  output         io_Pctrl_isclip_32,
  output         io_Pctrl_isClip,
  output         io_Pctrl_isSat_16,
  output         io_Pctrl_isSat_8,
  output         io_Pctrl_isSat_32,
  output         io_Pctrl_isSat_W,
  output         io_Pctrl_isSat,
  output         io_Pctrl_isCnt_16,
  output         io_Pctrl_isCnt_8,
  output         io_Pctrl_isCnt_32,
  output         io_Pctrl_isCnt,
  output         io_Pctrl_isSwap_16,
  output         io_Pctrl_isSwap_8,
  output         io_Pctrl_isSwap,
  output         io_Pctrl_isUnpack,
  output         io_Pctrl_isBitrev,
  output         io_Pctrl_isCmix,
  output         io_Pctrl_isInsertb,
  output         io_Pctrl_isPackbb,
  output         io_Pctrl_isPackbt,
  output         io_Pctrl_isPacktb,
  output         io_Pctrl_isPacktt,
  output         io_Pctrl_isPack,
  output [7:0]   io_Pctrl_isSub,
  output         io_Pctrl_isAdder,
  output         io_Pctrl_SrcSigned,
  output         io_Pctrl_Saturating,
  output         io_Pctrl_Translation,
  output         io_Pctrl_LessEqual,
  output         io_Pctrl_LessThan,
  output [79:0]  io_Pctrl_adderRes_ori,
  output [63:0]  io_Pctrl_adderRes,
  output [79:0]  io_Pctrl_adderRes_ori_drophighestbit,
  output         io_Pctrl_Round,
  output         io_Pctrl_ShiftSigned,
  output         io_Pctrl_Arithmetic,
  output         io_Pctrl_isMul_16,
  output         io_Pctrl_isMul_8,
  output         io_Pctrl_isMSW_3232,
  output         io_Pctrl_isMSW_3216,
  output         io_Pctrl_isS1632,
  output         io_Pctrl_isS1664,
  output         io_Pctrl_is832,
  output         io_Pctrl_is3264,
  output         io_Pctrl_is1664,
  output         io_Pctrl_isQ15orQ31,
  output         io_Pctrl_isC31,
  output         io_Pctrl_isQ15_64ONLY,
  output         io_Pctrl_isQ63_64ONLY,
  output         io_Pctrl_isMul_32_64ONLY,
  output         io_Pctrl_isPMA_64ONLY,
  output [17:0]  io_Pctrl_mulres9_0,
  output [17:0]  io_Pctrl_mulres9_1,
  output [17:0]  io_Pctrl_mulres9_2,
  output [17:0]  io_Pctrl_mulres9_3,
  output [33:0]  io_Pctrl_mulres17_0,
  output [33:0]  io_Pctrl_mulres17_1,
  output [65:0]  io_Pctrl_mulres33_0,
  output [129:0] io_Pctrl_mulres65_0
);
  wire [16:0] MulAdd17_0_io_in_srcs_0; // @[PIDU.scala 292:28]
  wire [16:0] MulAdd17_0_io_in_srcs_1; // @[PIDU.scala 292:28]
  wire [33:0] MulAdd17_0_io_out_result; // @[PIDU.scala 292:28]
  wire [16:0] MulAdd17_1_io_in_srcs_0; // @[PIDU.scala 293:28]
  wire [16:0] MulAdd17_1_io_in_srcs_1; // @[PIDU.scala 293:28]
  wire [33:0] MulAdd17_1_io_out_result; // @[PIDU.scala 293:28]
  wire [32:0] MulAdd33_0_io_in_srcs_0; // @[PIDU.scala 294:28]
  wire [32:0] MulAdd33_0_io_in_srcs_1; // @[PIDU.scala 294:28]
  wire [65:0] MulAdd33_0_io_out_result; // @[PIDU.scala 294:28]
  wire [64:0] MulAdd65_0_io_in_srcs_0; // @[PIDU.scala 295:28]
  wire [64:0] MulAdd65_0_io_in_srcs_1; // @[PIDU.scala 295:28]
  wire [129:0] MulAdd65_0_io_out_result; // @[PIDU.scala 295:28]
  wire [8:0] MulAdd9_0_io_in_srcs_0; // @[PIDU.scala 296:28]
  wire [8:0] MulAdd9_0_io_in_srcs_1; // @[PIDU.scala 296:28]
  wire [17:0] MulAdd9_0_io_out_result; // @[PIDU.scala 296:28]
  wire [8:0] MulAdd9_1_io_in_srcs_0; // @[PIDU.scala 297:28]
  wire [8:0] MulAdd9_1_io_in_srcs_1; // @[PIDU.scala 297:28]
  wire [17:0] MulAdd9_1_io_out_result; // @[PIDU.scala 297:28]
  wire [8:0] MulAdd9_2_io_in_srcs_0; // @[PIDU.scala 298:28]
  wire [8:0] MulAdd9_2_io_in_srcs_1; // @[PIDU.scala 298:28]
  wire [17:0] MulAdd9_2_io_out_result; // @[PIDU.scala 298:28]
  wire [8:0] MulAdd9_3_io_in_srcs_0; // @[PIDU.scala 299:28]
  wire [8:0] MulAdd9_3_io_in_srcs_1; // @[PIDU.scala 299:28]
  wire [17:0] MulAdd9_3_io_out_result; // @[PIDU.scala 299:28]
  wire  _T_1 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h2; // @[PIDU.scala 154:36]
  wire  _T_3 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h0; // @[PIDU.scala 154:61]
  wire  _T_5 = io_DecodeIn_ctrl_funct3 == 3'h1; // @[PIDU.scala 154:84]
  wire  _T_10 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0; // @[PIDU.scala 155:72]
  wire  _T_12 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4; // @[PIDU.scala 155:94]
  wire  _T_13 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4; // @[PIDU.scala 155:80]
  wire  _T_14 = _T_3 & (io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4); // @[PIDU.scala 155:51]
  wire  _T_15 = io_DecodeIn_ctrl_funct3 == 3'h2; // @[PIDU.scala 155:113]
  wire  _T_25 = io_DecodeIn_ctrl_funct3 == 3'h0; // @[PIDU.scala 156:113]
  wire  _T_28 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h4; // @[PIDU.scala 157:43]
  wire  _T_38 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h0; // @[PIDU.scala 158:36]
  wire  _T_40 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h2; // @[PIDU.scala 158:62]
  wire  _T_52 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h1; // @[PIDU.scala 160:36]
  wire  _T_71 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h1; // @[PIDU.scala 164:61]
  wire  _T_82 = _T_71 & _T_13; // @[PIDU.scala 165:51]
  wire  _T_96 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h5; // @[PIDU.scala 167:43]
  wire  _T_108 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h3; // @[PIDU.scala 168:62]
  wire  _T_133 = _T_40 & _T_13; // @[PIDU.scala 172:52]
  wire  _T_143 = _T_108 & _T_13; // @[PIDU.scala 173:52]
  wire  _T_166 = io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16; // @[PIDU.scala 176:41]
  wire  _T_170 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h3; // @[PIDU.scala 178:38]
  wire  _T_172 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h5; // @[PIDU.scala 178:63]
  wire  _T_173 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h3 | io_DecodeIn_ctrl_fuOpType[6:4] == 3'h5; // @[PIDU.scala 178:50]
  wire  _T_213 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h6; // @[PIDU.scala 184:44]
  wire  _T_223 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h7; // @[PIDU.scala 185:44]
  wire  _T_234 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h4; // @[PIDU.scala 188:40]
  wire  _T_236 = io_DecodeIn_ctrl_fuOpType[2:1] == 2'h0; // @[PIDU.scala 188:61]
  wire  _T_243 = io_DecodeIn_ctrl_fuOpType[2:1] == 2'h2; // @[PIDU.scala 189:61]
  wire  _T_255 = io_DecodeIn_cf_instr[6:0] == 7'h33; // @[PIDU.scala 190:130]
  wire  _T_258 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h9; // @[PIDU.scala 191:41]
  wire  _T_275 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h1; // @[PIDU.scala 196:35]
  wire  _T_277 = io_DecodeIn_ctrl_fuOpType[4:3] != 2'h0; // @[PIDU.scala 196:56]
  wire  _T_278 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h1 & io_DecodeIn_ctrl_fuOpType[4:3] != 2'h0; // @[PIDU.scala 196:43]
  wire  _T_295 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5; // @[PIDU.scala 198:35]
  wire  _T_297 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6; // @[PIDU.scala 198:56]
  wire  _T_298 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6; // @[PIDU.scala 198:43]
  wire  _T_301 = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6) & _T_108; // @[PIDU.scala 198:64]
  wire  _T_340 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h8; // @[PIDU.scala 202:81]
  wire  _T_341 = _T_278 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h8; // @[PIDU.scala 202:68]
  wire  _T_371 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h3; // @[PIDU.scala 205:35]
  wire  _T_385 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h2; // @[PIDU.scala 207:38]
  wire  _T_387 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hd; // @[PIDU.scala 207:64]
  wire  _T_390 = io_DecodeIn_ctrl_fuOpType[2:1] == 2'h1; // @[PIDU.scala 207:91]
  wire  _T_399 = io_DecodeIn_ctrl_funct3 == 3'h5; // @[PIDU.scala 209:76]
  wire  _T_431 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h7; // @[PIDU.scala 215:37]
  wire  _T_439 = io_DecodeIn_ctrl_fuOpType == 7'h56; // @[PIDU.scala 218:32]
  wire  _T_466 = io_DecodeIn_ctrl_fuOpType == 7'h57; // @[PIDU.scala 224:32]
  wire  _T_530 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'he & (_T_108 | _T_243) & _T_25; // @[PIDU.scala 235:105]
  wire  _T_556 = io_DecodeIn_ctrl_funct3 == 3'h4; // @[PIDU.scala 242:59]
  wire  _T_624 = io_DecodeIn_ctrl_fuOpType == 7'h27; // @[PIDU.scala 252:168]
  wire  _T_633 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hc; // @[PIDU.scala 254:37]
  wire  _T_635 = io_DecodeIn_ctrl_fuOpType[2:0] != 3'h7; // @[PIDU.scala 254:64]
  wire  _T_711 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h1; // @[PIDU.scala 261:72]
  wire  _T_747 = io_DecodeIn_ctrl_fuOpType[1:0] == 2'h1 | _T_258; // @[PIDU.scala 264:57]
  wire [15:0] _GEN_0 = _T_747 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 279:23 281:29]
  wire [15:0] _GEN_1 = _T_747 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 279:23 283:29]
  wire [15:0] _GEN_2 = _T_747 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 279:23 281:29]
  wire [15:0] _GEN_3 = _T_747 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 279:23 283:29]
  wire [63:0] _T_758 = {_GEN_3,_GEN_2,_GEN_1,_GEN_0}; // @[Cat.scala 30:58]
  wire  _T_760 = io_DecodeIn_ctrl_fuOpType[1:0] == 2'h3; // @[PIDU.scala 265:44]
  wire  _T_762 = io_DecodeIn_ctrl_fuOpType[6:3] != 4'hb; // @[PIDU.scala 263:44]
  wire [16:0] _T_765 = {io_DecodeIn_data_src1[15],io_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _T_766 = {1'h0,io_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_4 = _T_762 ? _T_765 : _T_766; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_771 = {io_DecodeIn_data_src1[31],io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _T_772 = {1'h0,io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_5 = _T_762 ? _T_771 : _T_772; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_778 = io_DecodeIn_data_src1[47] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_779 = {_T_778,io_DecodeIn_data_src1[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _T_780 = {17'h0,io_DecodeIn_data_src1[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_6 = _T_762 ? _T_779 : _T_780; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_786 = io_DecodeIn_data_src1[63] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_787 = {_T_786,io_DecodeIn_data_src1[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _T_788 = {49'h0,io_DecodeIn_data_src1[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_7 = _T_762 ? _T_787 : _T_788; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_793 = {_T_758[15],_T_758[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _T_794 = {1'h0,_T_758[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_8 = _T_762 ? _T_793 : _T_794; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_799 = {_T_758[31],_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _T_800 = {1'h0,_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_9 = _T_762 ? _T_799 : _T_800; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _T_806 = _T_758[47] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_807 = {_T_806,_T_758[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _T_808 = {17'h0,_T_758[47:32]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_10 = _T_762 ? _T_807 : _T_808; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_814 = _T_758[63] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_815 = {_T_814,_T_758[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _T_816 = {49'h0,_T_758[63:48]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_11 = _T_762 ? _T_815 : _T_816; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_856 = io_DecodeIn_data_src1[31] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_857 = {_T_856,io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _T_858 = {49'h0,io_DecodeIn_data_src1[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_17 = _T_762 ? _T_857 : _T_858; // @[PIDU.scala 268:24 269:15 271:15]
  wire [48:0] _T_870 = _T_758[31] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_871 = {_T_870,_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _T_872 = {49'h0,_T_758[31:16]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_19 = _T_762 ? _T_871 : _T_872; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _GEN_22 = _T_760 ? _GEN_4 : _GEN_4; // @[PIDU.scala 314:35 315:42 328:42]
  wire [16:0] _GEN_23 = _T_760 ? _GEN_5 : 17'h0; // @[PIDU.scala 302:22 314:35 316:42]
  wire [32:0] _GEN_24 = _T_760 ? _GEN_6 : 33'h0; // @[PIDU.scala 303:22 314:35 317:42]
  wire [64:0] _GEN_25 = _T_760 ? _GEN_7 : _GEN_17; // @[PIDU.scala 314:35 318:42 329:42]
  wire [16:0] _GEN_26 = _T_760 ? _GEN_8 : _GEN_8; // @[PIDU.scala 314:35 319:42 330:42]
  wire [16:0] _GEN_27 = _T_760 ? _GEN_9 : 17'h0; // @[PIDU.scala 302:22 314:35 320:42]
  wire [32:0] _GEN_28 = _T_760 ? _GEN_10 : 33'h0; // @[PIDU.scala 303:22 314:35 321:42]
  wire [64:0] _GEN_29 = _T_760 ? _GEN_11 : _GEN_19; // @[PIDU.scala 314:35 322:42 331:42]
  wire [7:0] _GEN_34 = _T_747 ? io_DecodeIn_data_src2[15:8] : io_DecodeIn_data_src2[7:0]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_35 = _T_747 ? io_DecodeIn_data_src2[7:0] : io_DecodeIn_data_src2[15:8]; // @[PIDU.scala 279:23 283:29]
  wire [7:0] _GEN_36 = _T_747 ? io_DecodeIn_data_src2[31:24] : io_DecodeIn_data_src2[23:16]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_37 = _T_747 ? io_DecodeIn_data_src2[23:16] : io_DecodeIn_data_src2[31:24]; // @[PIDU.scala 279:23 283:29]
  wire [7:0] _GEN_38 = _T_747 ? io_DecodeIn_data_src2[47:40] : io_DecodeIn_data_src2[39:32]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_39 = _T_747 ? io_DecodeIn_data_src2[39:32] : io_DecodeIn_data_src2[47:40]; // @[PIDU.scala 279:23 283:29]
  wire [7:0] _GEN_40 = _T_747 ? io_DecodeIn_data_src2[63:56] : io_DecodeIn_data_src2[55:48]; // @[PIDU.scala 279:23 281:29]
  wire [7:0] _GEN_41 = _T_747 ? io_DecodeIn_data_src2[55:48] : io_DecodeIn_data_src2[63:56]; // @[PIDU.scala 279:23 283:29]
  wire [63:0] _T_914 = {_GEN_41,_GEN_40,_GEN_39,_GEN_38,_GEN_37,_GEN_36,_GEN_35,_GEN_34}; // @[Cat.scala 30:58]
  wire [8:0] _T_921 = {io_DecodeIn_data_src1[7],io_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _T_922 = {1'h0,io_DecodeIn_data_src1[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_42 = _T_762 ? _T_921 : _T_922; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_927 = {io_DecodeIn_data_src1[15],io_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _T_928 = {1'h0,io_DecodeIn_data_src1[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_43 = _T_762 ? _T_927 : _T_928; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_933 = {io_DecodeIn_data_src1[23],io_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _T_934 = {1'h0,io_DecodeIn_data_src1[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_44 = _T_762 ? _T_933 : _T_934; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_939 = {io_DecodeIn_data_src1[31],io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _T_940 = {1'h0,io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_45 = _T_762 ? _T_939 : _T_940; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_946 = io_DecodeIn_data_src1[39] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_947 = {_T_946,io_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _T_948 = {9'h0,io_DecodeIn_data_src1[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_46 = _T_762 ? _T_947 : _T_948; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_954 = io_DecodeIn_data_src1[47] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_955 = {_T_954,io_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _T_956 = {9'h0,io_DecodeIn_data_src1[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_47 = _T_762 ? _T_955 : _T_956; // @[PIDU.scala 268:24 269:15 271:15]
  wire [24:0] _T_962 = io_DecodeIn_data_src1[55] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_963 = {_T_962,io_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _T_964 = {25'h0,io_DecodeIn_data_src1[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_48 = _T_762 ? _T_963 : _T_964; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_970 = io_DecodeIn_data_src1[63] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_971 = {_T_970,io_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _T_972 = {57'h0,io_DecodeIn_data_src1[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_49 = _T_762 ? _T_971 : _T_972; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_977 = {_T_914[7],_T_914[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _T_978 = {1'h0,_T_914[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_50 = _T_762 ? _T_977 : _T_978; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_983 = {_T_914[15],_T_914[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _T_984 = {1'h0,_T_914[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_51 = _T_762 ? _T_983 : _T_984; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_989 = {_T_914[23],_T_914[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _T_990 = {1'h0,_T_914[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_52 = _T_762 ? _T_989 : _T_990; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_995 = {_T_914[31],_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _T_996 = {1'h0,_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_53 = _T_762 ? _T_995 : _T_996; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1002 = _T_914[39] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1003 = {_T_1002,_T_914[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1004 = {9'h0,_T_914[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_54 = _T_762 ? _T_1003 : _T_1004; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1010 = _T_914[47] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1011 = {_T_1010,_T_914[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1012 = {9'h0,_T_914[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_55 = _T_762 ? _T_1011 : _T_1012; // @[PIDU.scala 268:24 269:15 271:15]
  wire [24:0] _T_1018 = _T_914[55] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1019 = {_T_1018,_T_914[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1020 = {25'h0,_T_914[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_56 = _T_762 ? _T_1019 : _T_1020; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1026 = _T_914[63] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1027 = {_T_1026,_T_914[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1028 = {57'h0,_T_914[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_57 = _T_762 ? _T_1027 : _T_1028; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1108 = io_DecodeIn_data_src1[31] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1109 = {_T_1108,io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1110 = {57'h0,io_DecodeIn_data_src1[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_69 = _T_762 ? _T_1109 : _T_1110; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1134 = _T_914[31] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1135 = {_T_1134,_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1136 = {57'h0,_T_914[31:24]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_73 = _T_762 ? _T_1135 : _T_1136; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_78 = _T_760 ? _GEN_42 : _GEN_42; // @[PIDU.scala 338:35 339:42 364:42]
  wire [8:0] _GEN_79 = _T_760 ? _GEN_43 : _GEN_43; // @[PIDU.scala 338:35 340:42 365:42]
  wire [8:0] _GEN_80 = _T_760 ? _GEN_44 : _GEN_44; // @[PIDU.scala 338:35 341:42 366:42]
  wire [8:0] _GEN_81 = _T_760 ? _GEN_45 : 9'h0; // @[PIDU.scala 308:22 338:35 342:42]
  wire [16:0] _GEN_82 = _T_760 ? _GEN_46 : 17'h0; // @[PIDU.scala 301:22 338:35 343:42]
  wire [16:0] _GEN_83 = _T_760 ? _GEN_47 : 17'h0; // @[PIDU.scala 302:22 338:35 344:42]
  wire [32:0] _GEN_84 = _T_760 ? _GEN_48 : 33'h0; // @[PIDU.scala 303:22 338:35 345:42]
  wire [64:0] _GEN_85 = _T_760 ? _GEN_49 : _GEN_69; // @[PIDU.scala 338:35 346:42 367:42]
  wire [8:0] _GEN_86 = _T_760 ? _GEN_50 : _GEN_50; // @[PIDU.scala 338:35 347:42 368:42]
  wire [8:0] _GEN_87 = _T_760 ? _GEN_51 : _GEN_51; // @[PIDU.scala 338:35 348:42 369:42]
  wire [8:0] _GEN_88 = _T_760 ? _GEN_52 : _GEN_52; // @[PIDU.scala 338:35 349:42 370:42]
  wire [8:0] _GEN_89 = _T_760 ? _GEN_53 : 9'h0; // @[PIDU.scala 308:22 338:35 350:42]
  wire [16:0] _GEN_90 = _T_760 ? _GEN_54 : 17'h0; // @[PIDU.scala 301:22 338:35 351:42]
  wire [16:0] _GEN_91 = _T_760 ? _GEN_55 : 17'h0; // @[PIDU.scala 302:22 338:35 352:42]
  wire [32:0] _GEN_92 = _T_760 ? _GEN_56 : 33'h0; // @[PIDU.scala 303:22 338:35 353:42]
  wire [64:0] _GEN_93 = _T_760 ? _GEN_57 : _GEN_73; // @[PIDU.scala 338:35 354:42 371:42]
  wire [32:0] _T_1172 = {io_DecodeIn_data_src1[31],io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1175 = {io_DecodeIn_data_src2[31],io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1181 = io_DecodeIn_data_src1[63] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1182 = {_T_1181,io_DecodeIn_data_src1[63:32]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1186 = io_DecodeIn_data_src2[63] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1187 = {_T_1186,io_DecodeIn_data_src2[63:32]}; // @[Cat.scala 30:58]
  wire  _T_1197 = _T_371 | _T_172 | _T_431; // @[PIDU.scala 388:81]
  wire [15:0] _T_1203 = _T_1197 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 390:52]
  wire [16:0] _T_1206 = _T_1203[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1207 = {_T_1206,_T_1203}; // @[Cat.scala 30:58]
  wire [15:0] _T_1217 = _T_1197 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 393:52]
  wire [48:0] _T_1220 = _T_1217[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1221 = {_T_1220,_T_1217}; // @[Cat.scala 30:58]
  wire  _T_1234 = io_DecodeIn_ctrl_fuOpType[6:3] < 4'h3 | _T_96 & _T_275 & _T_277; // @[PIDU.scala 396:44]
  wire  _T_1239 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h0 | _T_295; // @[PIDU.scala 398:50]
  wire  _T_1244 = _T_711 | _T_297; // @[PIDU.scala 399:50]
  wire [15:0] _T_1248 = _T_1244 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 400:55]
  wire [15:0] _T_1249 = _T_1239 ? io_DecodeIn_data_src1[15:0] : _T_1248; // @[PIDU.scala 400:37]
  wire [15:0] _T_1253 = _T_1244 ? io_DecodeIn_data_src1[47:32] : io_DecodeIn_data_src1[63:48]; // @[PIDU.scala 401:56]
  wire [15:0] _T_1254 = _T_1239 ? io_DecodeIn_data_src1[47:32] : _T_1253; // @[PIDU.scala 401:37]
  wire [15:0] _T_1257 = _T_1239 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 402:37]
  wire [15:0] _T_1260 = _T_1239 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 403:37]
  wire [16:0] _T_1263 = _T_1249[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1264 = {_T_1263,_T_1249}; // @[Cat.scala 30:58]
  wire [16:0] _T_1267 = _T_1257[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1268 = {_T_1267,_T_1257}; // @[Cat.scala 30:58]
  wire [48:0] _T_1273 = _T_1254[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1274 = {_T_1273,_T_1254}; // @[Cat.scala 30:58]
  wire [48:0] _T_1277 = _T_1260[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1278 = {_T_1277,_T_1260}; // @[Cat.scala 30:58]
  wire  _T_1288 = io_DecodeIn_ctrl_fuOpType == 7'h3e; // @[PIDU.scala 411:134]
  wire  _T_1289 = io_DecodeIn_ctrl_fuOpType == 7'h1d | io_DecodeIn_ctrl_fuOpType == 7'h25 | _T_624 |
    io_DecodeIn_ctrl_fuOpType == 7'h3c | io_DecodeIn_ctrl_fuOpType == 7'h3e; // @[PIDU.scala 411:126]
  wire [15:0] _T_1296 = _T_1289 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 413:71]
  wire [15:0] _T_1299 = _T_1289 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 413:105]
  wire [15:0] _T_1302 = _T_1289 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 413:139]
  wire [15:0] _T_1305 = _T_1289 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 413:174]
  wire [16:0] _T_1309 = {_T_1296[15],_T_1296}; // @[Cat.scala 30:58]
  wire [48:0] _T_1318 = _T_1299[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1319 = {_T_1318,_T_1299}; // @[Cat.scala 30:58]
  wire [16:0] _T_1328 = _T_1302[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1329 = {_T_1328,_T_1302}; // @[Cat.scala 30:58]
  wire [48:0] _T_1338 = _T_1305[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1339 = {_T_1338,_T_1305}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_102 = _T_1234 ? _T_1264 : _T_779; // @[PIDU.scala 397:27 404:42 420:42]
  wire [32:0] _GEN_103 = _T_1234 ? _T_1268 : _T_1329; // @[PIDU.scala 397:27 405:42 421:42]
  wire [64:0] _GEN_105 = _T_1234 ? _T_1274 : _T_787; // @[PIDU.scala 397:27 407:42 423:42]
  wire [64:0] _GEN_106 = _T_1234 ? _T_1278 : _T_1339; // @[PIDU.scala 397:27 408:42 424:42]
  wire [16:0] _GEN_108 = _T_1234 ? 17'h0 : _T_765; // @[PIDU.scala 301:22 397:27 414:42]
  wire [16:0] _GEN_109 = _T_1234 ? 17'h0 : _T_1309; // @[PIDU.scala 301:22 397:27 415:42]
  wire [64:0] _GEN_111 = _T_1234 ? 65'h0 : _T_857; // @[PIDU.scala 302:22 397:27 417:42]
  wire [64:0] _GEN_112 = _T_1234 ? 65'h0 : _T_1319; // @[PIDU.scala 302:22 397:27 418:42]
  wire [16:0] _T_1345 = io_DecodeIn_data_src2[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1346 = {_T_1345,io_DecodeIn_data_src2[15:0]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1350 = io_DecodeIn_data_src2[31] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1351 = {_T_1350,io_DecodeIn_data_src2[31:16]}; // @[Cat.scala 30:58]
  wire [48:0] _T_1357 = io_DecodeIn_data_src2[47] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1358 = {_T_1357,io_DecodeIn_data_src2[47:32]}; // @[Cat.scala 30:58]
  wire [48:0] _T_1362 = io_DecodeIn_data_src2[63] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1363 = {_T_1362,io_DecodeIn_data_src2[63:48]}; // @[Cat.scala 30:58]
  wire  _T_1370 = ~_T_213; // @[PIDU.scala 438:50]
  wire [8:0] _GEN_114 = _T_1370 ? _T_921 : _T_922; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_115 = _T_1370 ? _T_927 : _T_928; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_116 = _T_1370 ? _T_933 : _T_934; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _GEN_117 = _T_1370 ? _T_939 : _T_940; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _GEN_118 = _T_1370 ? _T_947 : _T_948; // @[PIDU.scala 268:24 269:15 271:15]
  wire [16:0] _GEN_119 = _T_1370 ? _T_955 : _T_956; // @[PIDU.scala 268:24 269:15 271:15]
  wire [32:0] _GEN_120 = _T_1370 ? _T_963 : _T_964; // @[PIDU.scala 268:24 269:15 271:15]
  wire [64:0] _GEN_121 = _T_1370 ? _T_971 : _T_972; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1420 = {io_DecodeIn_data_src2[7],io_DecodeIn_data_src2[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1421 = {1'h0,io_DecodeIn_data_src2[7:0]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_122 = _T_28 ? _T_1420 : _T_1421; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1424 = {io_DecodeIn_data_src2[15],io_DecodeIn_data_src2[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1425 = {1'h0,io_DecodeIn_data_src2[15:8]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_123 = _T_28 ? _T_1424 : _T_1425; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1428 = {io_DecodeIn_data_src2[23],io_DecodeIn_data_src2[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1429 = {1'h0,io_DecodeIn_data_src2[23:16]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_124 = _T_28 ? _T_1428 : _T_1429; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1432 = {io_DecodeIn_data_src2[31],io_DecodeIn_data_src2[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _T_1433 = {1'h0,io_DecodeIn_data_src2[31:24]}; // @[Cat.scala 30:58]
  wire [8:0] _GEN_125 = _T_28 ? _T_1432 : _T_1433; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1437 = io_DecodeIn_data_src2[39] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1438 = {_T_1437,io_DecodeIn_data_src2[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1439 = {9'h0,io_DecodeIn_data_src2[39:32]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_126 = _T_28 ? _T_1438 : _T_1439; // @[PIDU.scala 268:24 269:15 271:15]
  wire [8:0] _T_1443 = io_DecodeIn_data_src2[47] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [16:0] _T_1444 = {_T_1443,io_DecodeIn_data_src2[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _T_1445 = {9'h0,io_DecodeIn_data_src2[47:40]}; // @[Cat.scala 30:58]
  wire [16:0] _GEN_127 = _T_28 ? _T_1444 : _T_1445; // @[PIDU.scala 268:24 269:15 271:15]
  wire [24:0] _T_1449 = io_DecodeIn_data_src2[55] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1450 = {_T_1449,io_DecodeIn_data_src2[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _T_1451 = {25'h0,io_DecodeIn_data_src2[55:48]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_128 = _T_28 ? _T_1450 : _T_1451; // @[PIDU.scala 268:24 269:15 271:15]
  wire [56:0] _T_1455 = io_DecodeIn_data_src2[63] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1456 = {_T_1455,io_DecodeIn_data_src2[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1457 = {57'h0,io_DecodeIn_data_src2[63:56]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_129 = _T_28 ? _T_1456 : _T_1457; // @[PIDU.scala 268:24 269:15 271:15]
  wire  _T_1460 = ~io_DecodeIn_ctrl_fuOpType[4]; // @[PIDU.scala 464:30]
  wire [32:0] _T_1464 = {1'h0,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_130 = _T_1460 ? _T_1172 : _T_1464; // @[PIDU.scala 268:24 269:15 271:15]
  wire [64:0] _T_1470 = {33'h0,io_DecodeIn_data_src1[63:32]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_131 = _T_1460 ? _T_1182 : _T_1470; // @[PIDU.scala 268:24 269:15 271:15]
  wire [32:0] _T_1474 = {1'h0,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_132 = _T_1460 ? _T_1175 : _T_1474; // @[PIDU.scala 268:24 269:15 271:15]
  wire [64:0] _T_1480 = {33'h0,io_DecodeIn_data_src2[63:32]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_133 = _T_1460 ? _T_1187 : _T_1480; // @[PIDU.scala 268:24 269:15 271:15]
  wire  _T_1484 = io_DecodeIn_ctrl_fuOpType[4:3] == 2'h0; // @[PIDU.scala 474:36]
  wire  _T_1486 = io_DecodeIn_ctrl_fuOpType[4:3] == 2'h1; // @[PIDU.scala 475:36]
  wire [15:0] _T_1490 = _T_1486 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 476:55]
  wire [15:0] _T_1491 = _T_1484 ? io_DecodeIn_data_src1[15:0] : _T_1490; // @[PIDU.scala 476:37]
  wire [15:0] _T_1495 = _T_1486 ? io_DecodeIn_data_src1[47:32] : io_DecodeIn_data_src1[63:48]; // @[PIDU.scala 477:56]
  wire [15:0] _T_1496 = _T_1484 ? io_DecodeIn_data_src1[47:32] : _T_1495; // @[PIDU.scala 477:37]
  wire [15:0] _T_1499 = _T_1484 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 478:37]
  wire [15:0] _T_1502 = _T_1484 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 479:37]
  wire [16:0] _T_1505 = _T_1491[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1506 = {_T_1505,_T_1491}; // @[Cat.scala 30:58]
  wire [16:0] _T_1509 = _T_1499[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1510 = {_T_1509,_T_1499}; // @[Cat.scala 30:58]
  wire [48:0] _T_1515 = _T_1496[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1516 = {_T_1515,_T_1496}; // @[Cat.scala 30:58]
  wire [48:0] _T_1519 = _T_1502[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1520 = {_T_1519,_T_1502}; // @[Cat.scala 30:58]
  wire  _T_1527 = io_DecodeIn_ctrl_fuOpType == 7'h55 | io_DecodeIn_ctrl_fuOpType == 7'h4e | io_DecodeIn_ctrl_fuOpType
     == 7'h5e; // @[PIDU.scala 487:76]
  wire [15:0] _T_1534 = _T_1527 ? io_DecodeIn_data_src2[31:16] : io_DecodeIn_data_src2[15:0]; // @[PIDU.scala 489:71]
  wire [15:0] _T_1537 = _T_1527 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 489:105]
  wire [15:0] _T_1540 = _T_1527 ? io_DecodeIn_data_src2[63:48] : io_DecodeIn_data_src2[47:32]; // @[PIDU.scala 489:139]
  wire [15:0] _T_1543 = _T_1527 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 489:174]
  wire [16:0] _T_1547 = {_T_1534[15],_T_1534}; // @[Cat.scala 30:58]
  wire [48:0] _T_1556 = _T_1537[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1557 = {_T_1556,_T_1537}; // @[Cat.scala 30:58]
  wire [16:0] _T_1566 = _T_1540[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1567 = {_T_1566,_T_1540}; // @[Cat.scala 30:58]
  wire [48:0] _T_1576 = _T_1543[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1577 = {_T_1576,_T_1543}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_134 = _T_28 ? _T_1506 : _T_779; // @[PIDU.scala 473:27 480:42 496:42]
  wire [32:0] _GEN_135 = _T_28 ? _T_1510 : _T_1567; // @[PIDU.scala 473:27 481:42 497:42]
  wire [64:0] _GEN_137 = _T_28 ? _T_1516 : _T_787; // @[PIDU.scala 473:27 483:42 499:42]
  wire [64:0] _GEN_138 = _T_28 ? _T_1520 : _T_1577; // @[PIDU.scala 473:27 484:42 500:42]
  wire [16:0] _GEN_140 = _T_28 ? 17'h0 : _T_765; // @[PIDU.scala 301:22 473:27 490:42]
  wire [16:0] _GEN_141 = _T_28 ? 17'h0 : _T_1547; // @[PIDU.scala 301:22 473:27 491:42]
  wire [64:0] _GEN_143 = _T_28 ? 65'h0 : _T_857; // @[PIDU.scala 302:22 473:27 493:42]
  wire [64:0] _GEN_144 = _T_28 ? 65'h0 : _T_1557; // @[PIDU.scala 302:22 473:27 494:42]
  wire  _T_1586 = _T_71 ? _T_1486 : _T_1484; // @[PIDU.scala 505:25]
  wire  _T_1588 = io_DecodeIn_ctrl_fuOpType[4:3] == 2'h2; // @[PIDU.scala 506:48]
  wire  _T_1591 = _T_71 ? io_DecodeIn_ctrl_fuOpType[4:3] == 2'h2 : _T_1486; // @[PIDU.scala 506:25]
  wire [15:0] _T_1595 = _T_1591 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 507:51]
  wire [15:0] _T_1596 = _T_1586 ? io_DecodeIn_data_src1[15:0] : _T_1595; // @[PIDU.scala 507:33]
  wire [15:0] _T_1599 = _T_1586 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 508:33]
  wire [48:0] _T_1602 = _T_1596[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1603 = {_T_1602,_T_1596}; // @[Cat.scala 30:58]
  wire [48:0] _T_1606 = _T_1599[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1607 = {_T_1606,_T_1599}; // @[Cat.scala 30:58]
  wire  _T_1611 = io_DecodeIn_ctrl_fuOpType[6:3] != 4'hf; // @[PIDU.scala 513:59]
  wire [32:0] _T_1615 = io_DecodeIn_data_src1[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1616 = {_T_1615,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1617 = {33'h0,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_146 = _T_1611 ? _T_1616 : _T_1617; // @[PIDU.scala 268:24 269:15 271:15]
  wire [32:0] _T_1623 = io_DecodeIn_data_src2[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1624 = {_T_1623,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _T_1625 = {33'h0,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_147 = _T_1611 ? _T_1624 : _T_1625; // @[PIDU.scala 268:24 269:15 271:15]
  wire [15:0] _T_1635 = _T_1588 ? io_DecodeIn_data_src1[15:0] : io_DecodeIn_data_src1[31:16]; // @[PIDU.scala 519:51]
  wire [15:0] _T_1636 = _T_1486 ? io_DecodeIn_data_src1[15:0] : _T_1635; // @[PIDU.scala 519:33]
  wire [15:0] _T_1640 = _T_1588 ? io_DecodeIn_data_src1[47:32] : io_DecodeIn_data_src1[63:48]; // @[PIDU.scala 520:52]
  wire [15:0] _T_1641 = _T_1486 ? io_DecodeIn_data_src1[47:32] : _T_1640; // @[PIDU.scala 520:33]
  wire [15:0] _T_1644 = _T_1486 ? io_DecodeIn_data_src2[15:0] : io_DecodeIn_data_src2[31:16]; // @[PIDU.scala 521:33]
  wire [15:0] _T_1647 = _T_1486 ? io_DecodeIn_data_src2[47:32] : io_DecodeIn_data_src2[63:48]; // @[PIDU.scala 522:33]
  wire [16:0] _T_1650 = _T_1636[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1651 = {_T_1650,_T_1636}; // @[Cat.scala 30:58]
  wire [16:0] _T_1654 = _T_1644[15] ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12]
  wire [32:0] _T_1655 = {_T_1654,_T_1644}; // @[Cat.scala 30:58]
  wire [48:0] _T_1660 = _T_1641[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1661 = {_T_1660,_T_1641}; // @[Cat.scala 30:58]
  wire [48:0] _T_1664 = _T_1647[15] ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1665 = {_T_1664,_T_1647}; // @[Cat.scala 30:58]
  wire [31:0] _T_1672 = _T_1486 ? io_DecodeIn_data_src1[31:0] : io_DecodeIn_data_src1[63:32]; // @[PIDU.scala 531:32]
  wire [32:0] _T_1676 = _T_1672[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1677 = {_T_1676,_T_1672}; // @[Cat.scala 30:58]
  wire [31:0] _T_1691 = _T_1588 ? io_DecodeIn_data_src1[31:0] : io_DecodeIn_data_src1[63:32]; // @[PIDU.scala 539:50]
  wire [31:0] _T_1692 = _T_1486 ? io_DecodeIn_data_src1[31:0] : _T_1691; // @[PIDU.scala 539:32]
  wire [31:0] _T_1695 = _T_1486 ? io_DecodeIn_data_src2[31:0] : io_DecodeIn_data_src2[63:32]; // @[PIDU.scala 540:32]
  wire [32:0] _T_1698 = _T_1692[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1699 = {_T_1698,_T_1692}; // @[Cat.scala 30:58]
  wire [32:0] _T_1702 = _T_1695[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1703 = {_T_1702,_T_1695}; // @[Cat.scala 30:58]
  wire  _T_1712 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'h7; // @[PIDU.scala 545:87]
  wire  _T_1713 = _T_96 | _T_223 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h7; // @[PIDU.scala 545:74]
  wire [31:0] _T_1718 = _T_1713 ? io_DecodeIn_data_src2[63:32] : io_DecodeIn_data_src2[31:0]; // @[PIDU.scala 548:33]
  wire [31:0] _T_1721 = _T_1713 ? io_DecodeIn_data_src2[31:0] : io_DecodeIn_data_src2[63:32]; // @[PIDU.scala 549:33]
  wire [32:0] _T_1725 = {_T_1718[31],_T_1718}; // @[Cat.scala 30:58]
  wire [32:0] _T_1734 = _T_1721[31] ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _T_1735 = {_T_1734,_T_1721}; // @[Cat.scala 30:58]
  wire [32:0] _GEN_148 = io_Pctrl_isPMA_64ONLY ? _T_1172 : 33'h0; // @[PIDU.scala 303:22 544:42 550:38]
  wire [32:0] _GEN_149 = io_Pctrl_isPMA_64ONLY ? _T_1725 : 33'h0; // @[PIDU.scala 303:22 544:42 551:38]
  wire [64:0] _GEN_151 = io_Pctrl_isPMA_64ONLY ? _T_1182 : 65'h0; // @[PIDU.scala 304:22 544:42 553:38]
  wire [64:0] _GEN_152 = io_Pctrl_isPMA_64ONLY ? _T_1735 : 65'h0; // @[PIDU.scala 304:22 544:42 554:38]
  wire [64:0] _GEN_154 = io_Pctrl_isQ63_64ONLY ? _T_1699 : _GEN_151; // @[PIDU.scala 536:42 541:38]
  wire [64:0] _GEN_155 = io_Pctrl_isQ63_64ONLY ? _T_1703 : _GEN_152; // @[PIDU.scala 536:42 542:38]
  wire [32:0] _GEN_157 = io_Pctrl_isQ63_64ONLY ? 33'h0 : _GEN_148; // @[PIDU.scala 303:22 536:42]
  wire [32:0] _GEN_158 = io_Pctrl_isQ63_64ONLY ? 33'h0 : _GEN_149; // @[PIDU.scala 303:22 536:42]
  wire [64:0] _GEN_160 = io_Pctrl_isMul_32_64ONLY ? _T_1677 : _GEN_154; // @[PIDU.scala 529:45 533:38]
  wire [64:0] _GEN_161 = io_Pctrl_isMul_32_64ONLY ? _T_1187 : _GEN_155; // @[PIDU.scala 529:45 534:38]
  wire [32:0] _GEN_163 = io_Pctrl_isMul_32_64ONLY ? 33'h0 : _GEN_157; // @[PIDU.scala 303:22 529:45]
  wire [32:0] _GEN_164 = io_Pctrl_isMul_32_64ONLY ? 33'h0 : _GEN_158; // @[PIDU.scala 303:22 529:45]
  wire [32:0] _GEN_166 = io_Pctrl_isQ15_64ONLY ? _T_1651 : _GEN_163; // @[PIDU.scala 516:42 523:38]
  wire [32:0] _GEN_167 = io_Pctrl_isQ15_64ONLY ? _T_1655 : _GEN_164; // @[PIDU.scala 516:42 524:38]
  wire [64:0] _GEN_169 = io_Pctrl_isQ15_64ONLY ? _T_1661 : _GEN_160; // @[PIDU.scala 516:42 526:38]
  wire [64:0] _GEN_170 = io_Pctrl_isQ15_64ONLY ? _T_1665 : _GEN_161; // @[PIDU.scala 516:42 527:38]
  wire [64:0] _GEN_172 = io_Pctrl_isC31 ? _GEN_146 : _GEN_169; // @[PIDU.scala 512:35 513:38]
  wire [64:0] _GEN_173 = io_Pctrl_isC31 ? _GEN_147 : _GEN_170; // @[PIDU.scala 512:35 514:38]
  wire [32:0] _GEN_175 = io_Pctrl_isC31 ? 33'h0 : _GEN_166; // @[PIDU.scala 303:22 512:35]
  wire [32:0] _GEN_176 = io_Pctrl_isC31 ? 33'h0 : _GEN_167; // @[PIDU.scala 303:22 512:35]
  wire [64:0] _GEN_178 = io_Pctrl_isQ15orQ31 ? _T_1603 : _GEN_172; // @[PIDU.scala 503:40 509:38]
  wire [64:0] _GEN_179 = io_Pctrl_isQ15orQ31 ? _T_1607 : _GEN_173; // @[PIDU.scala 503:40 510:38]
  wire [32:0] _GEN_181 = io_Pctrl_isQ15orQ31 ? 33'h0 : _GEN_175; // @[PIDU.scala 303:22 503:40]
  wire [32:0] _GEN_182 = io_Pctrl_isQ15orQ31 ? 33'h0 : _GEN_176; // @[PIDU.scala 303:22 503:40]
  wire [32:0] _GEN_184 = io_Pctrl_is1664 ? _GEN_134 : _GEN_181; // @[PIDU.scala 471:36]
  wire [32:0] _GEN_185 = io_Pctrl_is1664 ? _GEN_135 : _GEN_182; // @[PIDU.scala 471:36]
  wire [64:0] _GEN_187 = io_Pctrl_is1664 ? _GEN_137 : _GEN_178; // @[PIDU.scala 471:36]
  wire [64:0] _GEN_188 = io_Pctrl_is1664 ? _GEN_138 : _GEN_179; // @[PIDU.scala 471:36]
  wire [16:0] _GEN_190 = io_Pctrl_is1664 ? _GEN_140 : 17'h0; // @[PIDU.scala 301:22 471:36]
  wire [16:0] _GEN_191 = io_Pctrl_is1664 ? _GEN_141 : 17'h0; // @[PIDU.scala 301:22 471:36]
  wire [64:0] _GEN_193 = io_Pctrl_is1664 ? _GEN_143 : 65'h0; // @[PIDU.scala 302:22 471:36]
  wire [64:0] _GEN_194 = io_Pctrl_is1664 ? _GEN_144 : 65'h0; // @[PIDU.scala 302:22 471:36]
  wire [32:0] _GEN_196 = io_Pctrl_is3264 ? _GEN_130 : _GEN_184; // @[PIDU.scala 462:36 465:38]
  wire [64:0] _GEN_197 = io_Pctrl_is3264 ? _GEN_131 : _GEN_187; // @[PIDU.scala 462:36 466:38]
  wire [32:0] _GEN_198 = io_Pctrl_is3264 ? _GEN_132 : _GEN_185; // @[PIDU.scala 462:36 467:38]
  wire [64:0] _GEN_199 = io_Pctrl_is3264 ? _GEN_133 : _GEN_188; // @[PIDU.scala 462:36 468:38]
  wire [16:0] _GEN_202 = io_Pctrl_is3264 ? 17'h0 : _GEN_190; // @[PIDU.scala 301:22 462:36]
  wire [16:0] _GEN_203 = io_Pctrl_is3264 ? 17'h0 : _GEN_191; // @[PIDU.scala 301:22 462:36]
  wire [64:0] _GEN_205 = io_Pctrl_is3264 ? 65'h0 : _GEN_193; // @[PIDU.scala 302:22 462:36]
  wire [64:0] _GEN_206 = io_Pctrl_is3264 ? 65'h0 : _GEN_194; // @[PIDU.scala 302:22 462:36]
  wire [8:0] _GEN_208 = io_Pctrl_is832 ? _GEN_114 : 9'h0; // @[PIDU.scala 305:22 434:35 438:38]
  wire [8:0] _GEN_209 = io_Pctrl_is832 ? _GEN_115 : 9'h0; // @[PIDU.scala 306:22 434:35 439:38]
  wire [8:0] _GEN_210 = io_Pctrl_is832 ? _GEN_116 : 9'h0; // @[PIDU.scala 307:22 434:35 440:38]
  wire [8:0] _GEN_211 = io_Pctrl_is832 ? _GEN_117 : 9'h0; // @[PIDU.scala 308:22 434:35 441:38]
  wire [16:0] _GEN_212 = io_Pctrl_is832 ? _GEN_118 : _GEN_202; // @[PIDU.scala 434:35 442:38]
  wire [64:0] _GEN_213 = io_Pctrl_is832 ? {{48'd0}, _GEN_119} : _GEN_205; // @[PIDU.scala 434:35 443:38]
  wire [32:0] _GEN_214 = io_Pctrl_is832 ? _GEN_120 : _GEN_196; // @[PIDU.scala 434:35 444:38]
  wire [64:0] _GEN_215 = io_Pctrl_is832 ? _GEN_121 : _GEN_197; // @[PIDU.scala 434:35 445:38]
  wire [8:0] _GEN_216 = io_Pctrl_is832 ? _GEN_122 : 9'h0; // @[PIDU.scala 305:22 434:35 446:38]
  wire [8:0] _GEN_217 = io_Pctrl_is832 ? _GEN_123 : 9'h0; // @[PIDU.scala 306:22 434:35 447:38]
  wire [8:0] _GEN_218 = io_Pctrl_is832 ? _GEN_124 : 9'h0; // @[PIDU.scala 307:22 434:35 448:38]
  wire [8:0] _GEN_219 = io_Pctrl_is832 ? _GEN_125 : 9'h0; // @[PIDU.scala 308:22 434:35 449:38]
  wire [16:0] _GEN_220 = io_Pctrl_is832 ? _GEN_126 : _GEN_203; // @[PIDU.scala 434:35 450:38]
  wire [64:0] _GEN_221 = io_Pctrl_is832 ? {{48'd0}, _GEN_127} : _GEN_206; // @[PIDU.scala 434:35 451:38]
  wire [32:0] _GEN_222 = io_Pctrl_is832 ? _GEN_128 : _GEN_198; // @[PIDU.scala 434:35 452:38]
  wire [64:0] _GEN_223 = io_Pctrl_is832 ? _GEN_129 : _GEN_199; // @[PIDU.scala 434:35 453:38]
  wire [32:0] _GEN_232 = io_Pctrl_isS1664 ? _T_1346 : _GEN_214; // @[PIDU.scala 427:37 428:38]
  wire [32:0] _GEN_233 = io_Pctrl_isS1664 ? _T_1351 : _GEN_222; // @[PIDU.scala 427:37 429:38]
  wire [64:0] _GEN_235 = io_Pctrl_isS1664 ? _T_1358 : _GEN_215; // @[PIDU.scala 427:37 431:38]
  wire [64:0] _GEN_236 = io_Pctrl_isS1664 ? _T_1363 : _GEN_223; // @[PIDU.scala 427:37 432:38]
  wire [8:0] _GEN_238 = io_Pctrl_isS1664 ? 9'h0 : _GEN_208; // @[PIDU.scala 305:22 427:37]
  wire [8:0] _GEN_239 = io_Pctrl_isS1664 ? 9'h0 : _GEN_209; // @[PIDU.scala 306:22 427:37]
  wire [8:0] _GEN_240 = io_Pctrl_isS1664 ? 9'h0 : _GEN_210; // @[PIDU.scala 307:22 427:37]
  wire [8:0] _GEN_241 = io_Pctrl_isS1664 ? 9'h0 : _GEN_211; // @[PIDU.scala 308:22 427:37]
  wire [16:0] _GEN_242 = io_Pctrl_isS1664 ? 17'h0 : _GEN_212; // @[PIDU.scala 301:22 427:37]
  wire [64:0] _GEN_243 = io_Pctrl_isS1664 ? 65'h0 : _GEN_213; // @[PIDU.scala 302:22 427:37]
  wire [8:0] _GEN_244 = io_Pctrl_isS1664 ? 9'h0 : _GEN_216; // @[PIDU.scala 305:22 427:37]
  wire [8:0] _GEN_245 = io_Pctrl_isS1664 ? 9'h0 : _GEN_217; // @[PIDU.scala 306:22 427:37]
  wire [8:0] _GEN_246 = io_Pctrl_isS1664 ? 9'h0 : _GEN_218; // @[PIDU.scala 307:22 427:37]
  wire [8:0] _GEN_247 = io_Pctrl_isS1664 ? 9'h0 : _GEN_219; // @[PIDU.scala 308:22 427:37]
  wire [16:0] _GEN_248 = io_Pctrl_isS1664 ? 17'h0 : _GEN_220; // @[PIDU.scala 301:22 427:37]
  wire [64:0] _GEN_249 = io_Pctrl_isS1664 ? 65'h0 : _GEN_221; // @[PIDU.scala 302:22 427:37]
  wire [32:0] _GEN_256 = io_Pctrl_isS1632 ? _GEN_102 : _GEN_232; // @[PIDU.scala 395:37]
  wire [32:0] _GEN_257 = io_Pctrl_isS1632 ? _GEN_103 : _GEN_233; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_259 = io_Pctrl_isS1632 ? _GEN_105 : _GEN_235; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_260 = io_Pctrl_isS1632 ? _GEN_106 : _GEN_236; // @[PIDU.scala 395:37]
  wire [16:0] _GEN_262 = io_Pctrl_isS1632 ? _GEN_108 : _GEN_242; // @[PIDU.scala 395:37]
  wire [16:0] _GEN_263 = io_Pctrl_isS1632 ? _GEN_109 : _GEN_248; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_265 = io_Pctrl_isS1632 ? _GEN_111 : _GEN_243; // @[PIDU.scala 395:37]
  wire [64:0] _GEN_266 = io_Pctrl_isS1632 ? _GEN_112 : _GEN_249; // @[PIDU.scala 395:37]
  wire [8:0] _GEN_268 = io_Pctrl_isS1632 ? 9'h0 : _GEN_238; // @[PIDU.scala 305:22 395:37]
  wire [8:0] _GEN_269 = io_Pctrl_isS1632 ? 9'h0 : _GEN_239; // @[PIDU.scala 306:22 395:37]
  wire [8:0] _GEN_270 = io_Pctrl_isS1632 ? 9'h0 : _GEN_240; // @[PIDU.scala 307:22 395:37]
  wire [8:0] _GEN_271 = io_Pctrl_isS1632 ? 9'h0 : _GEN_241; // @[PIDU.scala 308:22 395:37]
  wire [8:0] _GEN_272 = io_Pctrl_isS1632 ? 9'h0 : _GEN_244; // @[PIDU.scala 305:22 395:37]
  wire [8:0] _GEN_273 = io_Pctrl_isS1632 ? 9'h0 : _GEN_245; // @[PIDU.scala 306:22 395:37]
  wire [8:0] _GEN_274 = io_Pctrl_isS1632 ? 9'h0 : _GEN_246; // @[PIDU.scala 307:22 395:37]
  wire [8:0] _GEN_275 = io_Pctrl_isS1632 ? 9'h0 : _GEN_247; // @[PIDU.scala 308:22 395:37]
  wire [32:0] _GEN_280 = io_Pctrl_isMSW_3216 ? _T_1172 : _GEN_256; // @[PIDU.scala 386:40 389:38]
  wire [32:0] _GEN_281 = io_Pctrl_isMSW_3216 ? _T_1207 : _GEN_257; // @[PIDU.scala 386:40 390:38]
  wire [64:0] _GEN_283 = io_Pctrl_isMSW_3216 ? _T_1182 : _GEN_259; // @[PIDU.scala 386:40 392:38]
  wire [64:0] _GEN_284 = io_Pctrl_isMSW_3216 ? _T_1221 : _GEN_260; // @[PIDU.scala 386:40 393:38]
  wire [16:0] _GEN_286 = io_Pctrl_isMSW_3216 ? 17'h0 : _GEN_262; // @[PIDU.scala 301:22 386:40]
  wire [16:0] _GEN_287 = io_Pctrl_isMSW_3216 ? 17'h0 : _GEN_263; // @[PIDU.scala 301:22 386:40]
  wire [64:0] _GEN_289 = io_Pctrl_isMSW_3216 ? 65'h0 : _GEN_265; // @[PIDU.scala 302:22 386:40]
  wire [64:0] _GEN_290 = io_Pctrl_isMSW_3216 ? 65'h0 : _GEN_266; // @[PIDU.scala 302:22 386:40]
  wire [8:0] _GEN_292 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_268; // @[PIDU.scala 305:22 386:40]
  wire [8:0] _GEN_293 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_269; // @[PIDU.scala 306:22 386:40]
  wire [8:0] _GEN_294 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_270; // @[PIDU.scala 307:22 386:40]
  wire [8:0] _GEN_295 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_271; // @[PIDU.scala 308:22 386:40]
  wire [8:0] _GEN_296 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_272; // @[PIDU.scala 305:22 386:40]
  wire [8:0] _GEN_297 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_273; // @[PIDU.scala 306:22 386:40]
  wire [8:0] _GEN_298 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_274; // @[PIDU.scala 307:22 386:40]
  wire [8:0] _GEN_299 = io_Pctrl_isMSW_3216 ? 9'h0 : _GEN_275; // @[PIDU.scala 308:22 386:40]
  wire [32:0] _GEN_304 = io_Pctrl_isMSW_3232 ? _T_1172 : _GEN_280; // @[PIDU.scala 378:40 380:38]
  wire [32:0] _GEN_305 = io_Pctrl_isMSW_3232 ? _T_1175 : _GEN_281; // @[PIDU.scala 378:40 381:38]
  wire [64:0] _GEN_307 = io_Pctrl_isMSW_3232 ? _T_1182 : _GEN_283; // @[PIDU.scala 378:40 383:38]
  wire [64:0] _GEN_308 = io_Pctrl_isMSW_3232 ? _T_1187 : _GEN_284; // @[PIDU.scala 378:40 384:38]
  wire [16:0] _GEN_310 = io_Pctrl_isMSW_3232 ? 17'h0 : _GEN_286; // @[PIDU.scala 301:22 378:40]
  wire [16:0] _GEN_311 = io_Pctrl_isMSW_3232 ? 17'h0 : _GEN_287; // @[PIDU.scala 301:22 378:40]
  wire [64:0] _GEN_313 = io_Pctrl_isMSW_3232 ? 65'h0 : _GEN_289; // @[PIDU.scala 302:22 378:40]
  wire [64:0] _GEN_314 = io_Pctrl_isMSW_3232 ? 65'h0 : _GEN_290; // @[PIDU.scala 302:22 378:40]
  wire [8:0] _GEN_316 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_292; // @[PIDU.scala 305:22 378:40]
  wire [8:0] _GEN_317 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_293; // @[PIDU.scala 306:22 378:40]
  wire [8:0] _GEN_318 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_294; // @[PIDU.scala 307:22 378:40]
  wire [8:0] _GEN_319 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_295; // @[PIDU.scala 308:22 378:40]
  wire [8:0] _GEN_320 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_296; // @[PIDU.scala 305:22 378:40]
  wire [8:0] _GEN_321 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_297; // @[PIDU.scala 306:22 378:40]
  wire [8:0] _GEN_322 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_298; // @[PIDU.scala 307:22 378:40]
  wire [8:0] _GEN_323 = io_Pctrl_isMSW_3232 ? 9'h0 : _GEN_299; // @[PIDU.scala 308:22 378:40]
  wire [8:0] _GEN_328 = io_Pctrl_isMul_8 ? _GEN_78 : _GEN_316; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_329 = io_Pctrl_isMul_8 ? _GEN_79 : _GEN_317; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_330 = io_Pctrl_isMul_8 ? _GEN_80 : _GEN_318; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_331 = io_Pctrl_isMul_8 ? _GEN_81 : _GEN_319; // @[PIDU.scala 335:37]
  wire [16:0] _GEN_332 = io_Pctrl_isMul_8 ? _GEN_82 : _GEN_310; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_333 = io_Pctrl_isMul_8 ? {{48'd0}, _GEN_83} : _GEN_313; // @[PIDU.scala 335:37]
  wire [32:0] _GEN_334 = io_Pctrl_isMul_8 ? _GEN_84 : _GEN_304; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_335 = io_Pctrl_isMul_8 ? _GEN_85 : _GEN_307; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_336 = io_Pctrl_isMul_8 ? _GEN_86 : _GEN_320; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_337 = io_Pctrl_isMul_8 ? _GEN_87 : _GEN_321; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_338 = io_Pctrl_isMul_8 ? _GEN_88 : _GEN_322; // @[PIDU.scala 335:37]
  wire [8:0] _GEN_339 = io_Pctrl_isMul_8 ? _GEN_89 : _GEN_323; // @[PIDU.scala 335:37]
  wire [16:0] _GEN_340 = io_Pctrl_isMul_8 ? _GEN_90 : _GEN_311; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_341 = io_Pctrl_isMul_8 ? {{48'd0}, _GEN_91} : _GEN_314; // @[PIDU.scala 335:37]
  wire [32:0] _GEN_342 = io_Pctrl_isMul_8 ? _GEN_92 : _GEN_305; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_343 = io_Pctrl_isMul_8 ? _GEN_93 : _GEN_308; // @[PIDU.scala 335:37]
  wire [64:0] _GEN_353 = io_Pctrl_isMul_16 ? {{48'd0}, _GEN_23} : _GEN_333; // @[PIDU.scala 311:32]
  wire [64:0] _GEN_357 = io_Pctrl_isMul_16 ? {{48'd0}, _GEN_27} : _GEN_341; // @[PIDU.scala 311:32]
  wire  _T_1748 = io_Pctrl_isSub_64 | io_Pctrl_isSub_32 | io_Pctrl_isSub_16 | io_Pctrl_isSub_8 | io_Pctrl_isComp_16; // @[PIDU.scala 633:87]
  wire [1:0] _GEN_376 = io_Pctrl_isCrsa_32 | io_Pctrl_isStsa_32 ? 2'h2 : 2'h0; // @[PIDU.scala 632:20 642:56 643:23]
  wire [1:0] _GEN_377 = io_Pctrl_isCras_32 | io_Pctrl_isStas_32 ? 2'h1 : _GEN_376; // @[PIDU.scala 640:56 641:23]
  wire [3:0] _GEN_378 = io_Pctrl_isCrsa_16 | io_Pctrl_isStsa_16 ? 4'ha : {{2'd0}, _GEN_377}; // @[PIDU.scala 638:56 639:23]
  wire [3:0] _GEN_379 = io_Pctrl_isCras_16 | io_Pctrl_isStas_16 ? 4'h5 : _GEN_378; // @[PIDU.scala 636:56 637:23]
  wire  _T_1775 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hb; // @[PIDU.scala 648:104]
  wire  _T_1781 = ~io_Pctrl_isSt; // @[PIDU.scala 649:29]
  wire  _T_1787 = ~io_DecodeIn_ctrl_fuOpType[3]; // @[PIDU.scala 649:82]
  wire  _T_1804 = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8; // @[PIDU.scala 797:32]
  wire  _T_1811 = io_Pctrl_isPbs ? 1'h0 : io_Pctrl_SrcSigned; // @[PIDU.scala 798:74]
  wire  _T_1812 = io_Pctrl_isMaxMin_8 ? _T_1787 : _T_1811; // @[PIDU.scala 798:34]
  wire [8:0] _T_1817 = {{1'd0}, io_DecodeIn_data_src1[7:0]}; // @[PIDU.scala 671:57]
  wire  _GEN_384 = _T_1812 & _T_1817[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1831 = {{1'd0}, io_DecodeIn_data_src1[15:8]}; // @[PIDU.scala 671:57]
  wire  _GEN_388 = _T_1812 & _T_1831[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1845 = {{1'd0}, io_DecodeIn_data_src1[23:16]}; // @[PIDU.scala 671:57]
  wire  _GEN_392 = _T_1812 & _T_1845[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1859 = {{1'd0}, io_DecodeIn_data_src1[31:24]}; // @[PIDU.scala 671:57]
  wire  _GEN_396 = _T_1812 & _T_1859[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1873 = {{1'd0}, io_DecodeIn_data_src1[39:32]}; // @[PIDU.scala 671:57]
  wire  _GEN_400 = _T_1812 & _T_1873[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1887 = {{1'd0}, io_DecodeIn_data_src1[47:40]}; // @[PIDU.scala 671:57]
  wire  _GEN_404 = _T_1812 & _T_1887[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1901 = {{1'd0}, io_DecodeIn_data_src1[55:48]}; // @[PIDU.scala 671:57]
  wire  _GEN_408 = _T_1812 & _T_1901[7]; // @[PIDU.scala 673:28]
  wire [8:0] _T_1915 = {{1'd0}, io_DecodeIn_data_src1[63:56]}; // @[PIDU.scala 671:57]
  wire  _GEN_412 = _T_1812 & _T_1915[7]; // @[PIDU.scala 673:28]
  wire [30:0] _T_1933 = {1'h0,_GEN_412,_T_1915[7:0],1'h0,_GEN_408,_T_1901[7:0],1'h0,_GEN_404,_T_1887[7:0],1'h0}; // @[Cat.scala 30:58]
  wire [60:0] _T_1942 = {_T_1933,_GEN_400,_T_1873[7:0],1'h0,_GEN_396,_T_1859[7:0],1'h0,_GEN_392,_T_1845[7:0],1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_1947 = {_T_1942,_GEN_388,_T_1831[7:0],1'h0,_GEN_384,_T_1817[7:0]}; // @[Cat.scala 30:58]
  wire [7:0] _T_1952 = io_Pctrl_isSub[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1953 = io_DecodeIn_data_src2[7:0] ^ _T_1952; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_577 = {{7'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_1956 = _T_1953 + _GEN_577; // @[PIDU.scala 671:57]
  wire  _T_1962 = io_Pctrl_isSub[0] & _T_1956 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_414 = io_Pctrl_isSub[0] & _T_1956 == 8'h80 ? 1'h0 : _T_1956[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_1965 = io_Pctrl_isSub[0] & _T_1956 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_416 = _T_1812 ? _GEN_414 : _T_1965; // @[PIDU.scala 673:28]
  wire [7:0] _T_1971 = io_Pctrl_isSub[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1972 = io_DecodeIn_data_src2[15:8] ^ _T_1971; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_578 = {{7'd0}, io_Pctrl_isSub[1]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_1975 = _T_1972 + _GEN_578; // @[PIDU.scala 671:57]
  wire  _T_1981 = io_Pctrl_isSub[1] & _T_1975 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_418 = io_Pctrl_isSub[1] & _T_1975 == 8'h80 ? 1'h0 : _T_1975[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_1984 = io_Pctrl_isSub[1] & _T_1975 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_420 = _T_1812 ? _GEN_418 : _T_1984; // @[PIDU.scala 673:28]
  wire [7:0] _T_1990 = io_Pctrl_isSub[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1991 = io_DecodeIn_data_src2[23:16] ^ _T_1990; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_579 = {{7'd0}, io_Pctrl_isSub[2]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_1994 = _T_1991 + _GEN_579; // @[PIDU.scala 671:57]
  wire  _T_2000 = io_Pctrl_isSub[2] & _T_1994 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_422 = io_Pctrl_isSub[2] & _T_1994 == 8'h80 ? 1'h0 : _T_1994[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2003 = io_Pctrl_isSub[2] & _T_1994 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_424 = _T_1812 ? _GEN_422 : _T_2003; // @[PIDU.scala 673:28]
  wire [7:0] _T_2009 = io_Pctrl_isSub[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2010 = io_DecodeIn_data_src2[31:24] ^ _T_2009; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_580 = {{7'd0}, io_Pctrl_isSub[3]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2013 = _T_2010 + _GEN_580; // @[PIDU.scala 671:57]
  wire  _T_2019 = io_Pctrl_isSub[3] & _T_2013 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_426 = io_Pctrl_isSub[3] & _T_2013 == 8'h80 ? 1'h0 : _T_2013[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2022 = io_Pctrl_isSub[3] & _T_2013 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_428 = _T_1812 ? _GEN_426 : _T_2022; // @[PIDU.scala 673:28]
  wire [7:0] _T_2028 = io_Pctrl_isSub[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2029 = io_DecodeIn_data_src2[39:32] ^ _T_2028; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_581 = {{7'd0}, io_Pctrl_isSub[4]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2032 = _T_2029 + _GEN_581; // @[PIDU.scala 671:57]
  wire  _T_2038 = io_Pctrl_isSub[4] & _T_2032 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_430 = io_Pctrl_isSub[4] & _T_2032 == 8'h80 ? 1'h0 : _T_2032[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2041 = io_Pctrl_isSub[4] & _T_2032 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_432 = _T_1812 ? _GEN_430 : _T_2041; // @[PIDU.scala 673:28]
  wire [7:0] _T_2047 = io_Pctrl_isSub[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2048 = io_DecodeIn_data_src2[47:40] ^ _T_2047; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_582 = {{7'd0}, io_Pctrl_isSub[5]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2051 = _T_2048 + _GEN_582; // @[PIDU.scala 671:57]
  wire  _T_2057 = io_Pctrl_isSub[5] & _T_2051 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_434 = io_Pctrl_isSub[5] & _T_2051 == 8'h80 ? 1'h0 : _T_2051[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2060 = io_Pctrl_isSub[5] & _T_2051 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_436 = _T_1812 ? _GEN_434 : _T_2060; // @[PIDU.scala 673:28]
  wire [7:0] _T_2066 = io_Pctrl_isSub[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2067 = io_DecodeIn_data_src2[55:48] ^ _T_2066; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_583 = {{7'd0}, io_Pctrl_isSub[6]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2070 = _T_2067 + _GEN_583; // @[PIDU.scala 671:57]
  wire  _T_2076 = io_Pctrl_isSub[6] & _T_2070 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_438 = io_Pctrl_isSub[6] & _T_2070 == 8'h80 ? 1'h0 : _T_2070[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2079 = io_Pctrl_isSub[6] & _T_2070 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_440 = _T_1812 ? _GEN_438 : _T_2079; // @[PIDU.scala 673:28]
  wire [7:0] _T_2085 = io_Pctrl_isSub[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_2086 = io_DecodeIn_data_src2[63:56] ^ _T_2085; // @[PIDU.scala 671:32]
  wire [7:0] _GEN_584 = {{7'd0}, io_Pctrl_isSub[7]}; // @[PIDU.scala 671:57]
  wire [7:0] _T_2089 = _T_2086 + _GEN_584; // @[PIDU.scala 671:57]
  wire  _T_2095 = io_Pctrl_isSub[7] & _T_2089 == 8'h80; // @[PIDU.scala 675:31]
  wire  _GEN_442 = io_Pctrl_isSub[7] & _T_2089 == 8'h80 ? 1'h0 : _T_2089[7]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2098 = io_Pctrl_isSub[7] & _T_2089 != 8'h0; // @[PIDU.scala 678:31]
  wire  _GEN_444 = _T_1812 ? _GEN_442 : _T_2098; // @[PIDU.scala 673:28]
  wire [30:0] _T_2108 = {1'h0,_GEN_444,_T_2089,1'h0,_GEN_440,_T_2070,1'h0,_GEN_436,_T_2051,1'h0}; // @[Cat.scala 30:58]
  wire [60:0] _T_2117 = {_T_2108,_GEN_432,_T_2032,1'h0,_GEN_428,_T_2013,1'h0,_GEN_424,_T_1994,1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_2122 = {_T_2117,_GEN_420,_T_1975,1'h0,_GEN_416,_T_1956}; // @[Cat.scala 30:58]
  wire [29:0] _T_2221 = {3'h0,_T_1915[6:0],1'h0,1'h0,1'h0,_T_1901[6:0],1'h0,1'h0,1'h0,_T_1887[6:0]}; // @[Cat.scala 30:58]
  wire [50:0] _T_2230 = {_T_2221,1'h0,1'h0,1'h0,_T_1873[6:0],1'h0,1'h0,1'h0,_T_1859[6:0],1'h0}; // @[Cat.scala 30:58]
  wire [71:0] _T_2239 = {_T_2230,1'h0,1'h0,_T_1845[6:0],1'h0,1'h0,1'h0,_T_1831[6:0],1'h0,1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_2241 = {_T_2239,1'h0,_T_1817[6:0]}; // @[Cat.scala 30:58]
  wire [22:0] _T_2371 = {2'h0,_T_2095,_T_2089[6:0],1'h0,1'h0,_T_2076,_T_2070[6:0],1'h0,1'h0,_T_2057}; // @[Cat.scala 30:58]
  wire [49:0] _T_2380 = {_T_2371,_T_2051[6:0],1'h0,1'h0,_T_2038,_T_2032[6:0],1'h0,1'h0,_T_2019,_T_2013[6:0]}; // @[Cat.scala 30:58]
  wire [70:0] _T_2389 = {_T_2380,1'h0,1'h0,_T_2000,_T_1994[6:0],1'h0,1'h0,_T_1981,_T_1975[6:0],1'h0}; // @[Cat.scala 30:58]
  wire [79:0] _T_2392 = {_T_2389,1'h0,_T_1962,_T_1956[6:0]}; // @[Cat.scala 30:58]
  wire  _T_2395 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16; // @[PIDU.scala 803:81]
  wire  _T_2402 = io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15; // @[PIDU.scala 804:51]
  wire [63:0] _T_2405 = {48'h0,io_DecodeIn_data_src1[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2406 = io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15 ? _T_2405 : io_DecodeIn_data_src1; // @[PIDU.scala 804:31]
  wire [63:0] _T_2410 = {48'h0,io_DecodeIn_data_src2[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2411 = _T_2402 ? _T_2410 : io_DecodeIn_data_src2; // @[PIDU.scala 805:31]
  wire  _T_2417 = io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15 ? _T_1787 : io_Pctrl_SrcSigned; // @[PIDU.scala 806:34]
  wire [16:0] _T_2424 = {{1'd0}, _T_2406[15:0]}; // @[PIDU.scala 671:57]
  wire  _GEN_480 = _T_2417 & _T_2424[15]; // @[PIDU.scala 673:28]
  wire [16:0] _T_2438 = {{1'd0}, _T_2406[31:16]}; // @[PIDU.scala 671:57]
  wire  _GEN_484 = _T_2417 & _T_2438[15]; // @[PIDU.scala 673:28]
  wire [16:0] _T_2452 = {{1'd0}, _T_2406[47:32]}; // @[PIDU.scala 671:57]
  wire  _GEN_488 = _T_2417 & _T_2452[15]; // @[PIDU.scala 673:28]
  wire [16:0] _T_2466 = {{1'd0}, _T_2406[63:48]}; // @[PIDU.scala 671:57]
  wire  _GEN_492 = _T_2417 & _T_2466[15]; // @[PIDU.scala 673:28]
  wire [54:0] _T_2484 = {1'h0,_GEN_492,_T_2466[15:0],1'h0,_GEN_488,_T_2452[15:0],1'h0,_GEN_484,_T_2438[15:0],1'h0}; // @[Cat.scala 30:58]
  wire [71:0] _T_2486 = {_T_2484,_GEN_480,_T_2424[15:0]}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_493 = _T_166 ? _T_2411[31:16] : _T_2411[15:0]; // @[PIDU.scala 663:21 664:23 666:29]
  wire [15:0] _T_2491 = io_Pctrl_isSub[0] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2492 = _GEN_493 ^ _T_2491; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_593 = {{15'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2495 = _T_2492 + _GEN_593; // @[PIDU.scala 671:57]
  wire  _T_2501 = io_Pctrl_isSub[0] & _T_2495 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_494 = io_Pctrl_isSub[0] & _T_2495 == 16'h8000 ? 1'h0 : _T_2495[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2504 = io_Pctrl_isSub[0] & _T_2495 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_496 = _T_2417 ? _GEN_494 : _T_2504; // @[PIDU.scala 673:28]
  wire [15:0] _GEN_497 = _T_166 ? _T_2411[15:0] : _T_2411[31:16]; // @[PIDU.scala 663:21 664:23 668:29]
  wire [15:0] _T_2510 = io_Pctrl_isSub[1] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2511 = _GEN_497 ^ _T_2510; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_594 = {{15'd0}, io_Pctrl_isSub[1]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2514 = _T_2511 + _GEN_594; // @[PIDU.scala 671:57]
  wire  _T_2520 = io_Pctrl_isSub[1] & _T_2514 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_498 = io_Pctrl_isSub[1] & _T_2514 == 16'h8000 ? 1'h0 : _T_2514[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2523 = io_Pctrl_isSub[1] & _T_2514 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_500 = _T_2417 ? _GEN_498 : _T_2523; // @[PIDU.scala 673:28]
  wire [15:0] _GEN_501 = _T_166 ? _T_2411[63:48] : _T_2411[47:32]; // @[PIDU.scala 663:21 664:23 666:29]
  wire [15:0] _T_2529 = io_Pctrl_isSub[2] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2530 = _GEN_501 ^ _T_2529; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_595 = {{15'd0}, io_Pctrl_isSub[2]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2533 = _T_2530 + _GEN_595; // @[PIDU.scala 671:57]
  wire  _T_2539 = io_Pctrl_isSub[2] & _T_2533 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_502 = io_Pctrl_isSub[2] & _T_2533 == 16'h8000 ? 1'h0 : _T_2533[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2542 = io_Pctrl_isSub[2] & _T_2533 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_504 = _T_2417 ? _GEN_502 : _T_2542; // @[PIDU.scala 673:28]
  wire [15:0] _GEN_505 = _T_166 ? _T_2411[47:32] : _T_2411[63:48]; // @[PIDU.scala 663:21 664:23 668:29]
  wire [15:0] _T_2548 = io_Pctrl_isSub[3] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_2549 = _GEN_505 ^ _T_2548; // @[PIDU.scala 671:32]
  wire [15:0] _GEN_596 = {{15'd0}, io_Pctrl_isSub[3]}; // @[PIDU.scala 671:57]
  wire [15:0] _T_2552 = _T_2549 + _GEN_596; // @[PIDU.scala 671:57]
  wire  _T_2558 = io_Pctrl_isSub[3] & _T_2552 == 16'h8000; // @[PIDU.scala 675:31]
  wire  _GEN_506 = io_Pctrl_isSub[3] & _T_2552 == 16'h8000 ? 1'h0 : _T_2552[15]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2561 = io_Pctrl_isSub[3] & _T_2552 != 16'h0; // @[PIDU.scala 678:31]
  wire  _GEN_508 = _T_2417 ? _GEN_506 : _T_2561; // @[PIDU.scala 673:28]
  wire [54:0] _T_2571 = {1'h0,_GEN_508,_T_2552,1'h0,_GEN_504,_T_2533,1'h0,_GEN_500,_T_2514,1'h0}; // @[Cat.scala 30:58]
  wire [71:0] _T_2573 = {_T_2571,_GEN_496,_T_2495}; // @[Cat.scala 30:58]
  wire [53:0] _T_2628 = {3'h0,_T_2466[14:0],1'h0,1'h0,1'h0,_T_2452[14:0],1'h0,1'h0,1'h0,_T_2438[14:0]}; // @[Cat.scala 30:58]
  wire [71:0] _T_2632 = {_T_2628,1'h0,1'h0,1'h0,_T_2424[14:0]}; // @[Cat.scala 30:58]
  wire [38:0] _T_2702 = {2'h0,_T_2558,_T_2552[14:0],1'h0,1'h0,_T_2539,_T_2533[14:0],1'h0,1'h0,_T_2520}; // @[Cat.scala 30:58]
  wire [71:0] _T_2707 = {_T_2702,_T_2514[14:0],1'h0,1'h0,_T_2501,_T_2495[14:0]}; // @[Cat.scala 30:58]
  wire  _T_2710 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32; // @[PIDU.scala 812:81]
  wire  _T_2720 = io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31; // @[PIDU.scala 813:93]
  wire [63:0] _T_2723 = {32'h0,io_DecodeIn_data_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2724 = io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2723 :
    io_DecodeIn_data_src1; // @[PIDU.scala 813:31]
  wire [63:0] _T_2730 = {32'h0,io_DecodeIn_data_src2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2731 = _T_2720 ? _T_2730 : io_DecodeIn_data_src2; // @[PIDU.scala 814:31]
  wire  _T_2740 = io_Pctrl_isMaxMin_32 ? io_DecodeIn_ctrl_fuOpType[3] : io_Pctrl_SrcSigned; // @[PIDU.scala 815:135]
  wire  _T_2741 = _T_2720 ? _T_1787 : _T_2740; // @[PIDU.scala 815:34]
  wire  _T_2742 = io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32; // @[PIDU.scala 816:50]
  wire [32:0] _T_2748 = {{1'd0}, _T_2724[31:0]}; // @[PIDU.scala 671:57]
  wire  _GEN_528 = _T_2741 & _T_2748[31]; // @[PIDU.scala 673:28]
  wire [32:0] _T_2762 = {{1'd0}, _T_2724[63:32]}; // @[PIDU.scala 671:57]
  wire  _GEN_532 = _T_2741 & _T_2762[31]; // @[PIDU.scala 673:28]
  wire [67:0] _T_2776 = {1'h0,_GEN_532,_T_2762[31:0],1'h0,_GEN_528,_T_2748[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_533 = _T_2742 ? _T_2731[63:32] : _T_2731[31:0]; // @[PIDU.scala 663:21 664:23 666:29]
  wire [31:0] _T_2781 = io_Pctrl_isSub[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2782 = _GEN_533 ^ _T_2781; // @[PIDU.scala 671:32]
  wire [31:0] _GEN_601 = {{31'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [31:0] _T_2785 = _T_2782 + _GEN_601; // @[PIDU.scala 671:57]
  wire  _T_2791 = io_Pctrl_isSub[0] & _T_2785 == 32'h80000000; // @[PIDU.scala 675:31]
  wire  _GEN_534 = io_Pctrl_isSub[0] & _T_2785 == 32'h80000000 ? 1'h0 : _T_2785[31]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2794 = io_Pctrl_isSub[0] & _T_2785 != 32'h0; // @[PIDU.scala 678:31]
  wire  _GEN_536 = _T_2741 ? _GEN_534 : _T_2794; // @[PIDU.scala 673:28]
  wire [31:0] _GEN_537 = _T_2742 ? _T_2731[31:0] : _T_2731[63:32]; // @[PIDU.scala 663:21 664:23 668:29]
  wire [31:0] _T_2800 = io_Pctrl_isSub[1] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2801 = _GEN_537 ^ _T_2800; // @[PIDU.scala 671:32]
  wire [31:0] _GEN_602 = {{31'd0}, io_Pctrl_isSub[1]}; // @[PIDU.scala 671:57]
  wire [31:0] _T_2804 = _T_2801 + _GEN_602; // @[PIDU.scala 671:57]
  wire  _T_2810 = io_Pctrl_isSub[1] & _T_2804 == 32'h80000000; // @[PIDU.scala 675:31]
  wire  _GEN_538 = io_Pctrl_isSub[1] & _T_2804 == 32'h80000000 ? 1'h0 : _T_2804[31]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2813 = io_Pctrl_isSub[1] & _T_2804 != 32'h0; // @[PIDU.scala 678:31]
  wire  _GEN_540 = _T_2741 ? _GEN_538 : _T_2813; // @[PIDU.scala 673:28]
  wire [67:0] _T_2819 = {1'h0,_GEN_540,_T_2804,1'h0,_GEN_536,_T_2785}; // @[Cat.scala 30:58]
  wire [67:0] _T_2848 = {3'h0,_T_2762[30:0],1'h0,1'h0,1'h0,_T_2748[30:0]}; // @[Cat.scala 30:58]
  wire [67:0] _T_2885 = {2'h0,_T_2810,_T_2804[30:0],1'h0,1'h0,_T_2791,_T_2785[30:0]}; // @[Cat.scala 30:58]
  wire  _T_2889 = io_Pctrl_isMaxMin_XLEN | io_Pctrl_isAve | io_Pctrl_SrcSigned; // @[PIDU.scala 822:34]
  wire [64:0] _T_2893 = {{1'd0}, io_DecodeIn_data_src1}; // @[PIDU.scala 671:57]
  wire  _GEN_551 = _T_2889 & _T_2893[63]; // @[PIDU.scala 673:28]
  wire [65:0] _T_2904 = {1'h0,_GEN_551,_T_2893[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2908 = io_Pctrl_isSub[0] ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2909 = io_DecodeIn_data_src2 ^ _T_2908; // @[PIDU.scala 671:32]
  wire [63:0] _GEN_605 = {{63'd0}, io_Pctrl_isSub[0]}; // @[PIDU.scala 671:57]
  wire [63:0] _T_2912 = _T_2909 + _GEN_605; // @[PIDU.scala 671:57]
  wire  _T_2918 = io_Pctrl_isSub[0] & _T_2912 == 64'h8000000000000000; // @[PIDU.scala 675:31]
  wire  _GEN_552 = io_Pctrl_isSub[0] & _T_2912 == 64'h8000000000000000 ? 1'h0 : _T_2912[63]; // @[PIDU.scala 674:27 675:{71,82}]
  wire  _T_2921 = io_Pctrl_isSub[0] & _T_2912 != 64'h0; // @[PIDU.scala 678:31]
  wire  _GEN_554 = _T_2889 ? _GEN_552 : _T_2921; // @[PIDU.scala 673:28]
  wire [65:0] _T_2924 = {1'h0,_GEN_554,_T_2912}; // @[Cat.scala 30:58]
  wire [65:0] _T_2937 = {3'h0,_T_2893[62:0]}; // @[Cat.scala 30:58]
  wire [65:0] _T_2954 = {2'h0,_T_2918,_T_2912[62:0]}; // @[Cat.scala 30:58]
  wire [67:0] _GEN_561 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2776 : {{2'd0}, _T_2904}; // @[PIDU.scala 812:251 817:18]
  wire [67:0] _GEN_562 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2819 : {{2'd0}, _T_2924}; // @[PIDU.scala 812:251 818:18]
  wire [67:0] _GEN_563 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2848 : {{2'd0}, _T_2937}; // @[PIDU.scala 812:251 819:33]
  wire [67:0] _GEN_564 = io_Pctrl_isAdd_32 | io_Pctrl_isSub_32 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32 |
    io_Pctrl_isStas_32 | io_Pctrl_isStsa_32 | io_Pctrl_isMaxMin_32 | io_Pctrl_isAdd_Q31 | io_Pctrl_isSub_Q31 |
    io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 ? _T_2885 : {{2'd0}, _T_2954}; // @[PIDU.scala 812:251 820:33]
  wire [71:0] _GEN_565 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2486 : {{4'd0}, _GEN_561}; // @[PIDU.scala 803:231 808:18]
  wire [71:0] _GEN_566 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2573 : {{4'd0}, _GEN_562}; // @[PIDU.scala 803:231 809:18]
  wire [71:0] _GEN_567 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2632 : {{4'd0}, _GEN_563}; // @[PIDU.scala 803:231 810:33]
  wire [71:0] _GEN_568 = io_Pctrl_isAdd_16 | io_Pctrl_isSub_16 | io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 |
    io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isComp_16 | io_Pctrl_isMaxMin_16 | io_Pctrl_isAdd_Q15 |
    io_Pctrl_isSub_Q15 ? _T_2707 : {{4'd0}, _GEN_564}; // @[PIDU.scala 803:231 811:33]
  wire [79:0] add1 = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 | io_Pctrl_isPbs ?
    _T_1947 : {{8'd0}, _GEN_565}; // @[PIDU.scala 797:111 799:18]
  wire [79:0] add2 = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 | io_Pctrl_isPbs ?
    _T_2122 : {{8'd0}, _GEN_566}; // @[PIDU.scala 797:111 800:18]
  wire [79:0] add1_drophighestbit = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 |
    io_Pctrl_isPbs ? _T_2241 : {{8'd0}, _GEN_567}; // @[PIDU.scala 797:111 801:33]
  wire [79:0] add2_drophighestbit = io_Pctrl_isAdd_8 | io_Pctrl_isSub_8 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin_8 |
    io_Pctrl_isPbs ? _T_2392 : {{8'd0}, _GEN_568}; // @[PIDU.scala 797:111 802:33]
  wire [80:0] _T_2955 = add1 + add2; // @[PIDU.scala 840:35]
  wire [80:0] _T_2956 = add1_drophighestbit + add2_drophighestbit; // @[PIDU.scala 841:65]
  wire [63:0] _T_2973 = {io_Pctrl_adderRes_ori[77:70],io_Pctrl_adderRes_ori[67:60],io_Pctrl_adderRes_ori[57:50],
    io_Pctrl_adderRes_ori[47:40],io_Pctrl_adderRes_ori[37:30],io_Pctrl_adderRes_ori[27:20],io_Pctrl_adderRes_ori[17:10],
    io_Pctrl_adderRes_ori[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_2987 = {io_Pctrl_adderRes_ori[69:54],io_Pctrl_adderRes_ori[51:36],io_Pctrl_adderRes_ori[33:18],
    io_Pctrl_adderRes_ori[15:0]}; // @[Cat.scala 30:58]
  wire  _T_2991 = _T_2710 | io_Pctrl_isAdd_Q31; // @[PIDU.scala 862:98]
  wire [63:0] _T_2999 = {io_Pctrl_adderRes_ori[65:34],io_Pctrl_adderRes_ori[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_574 = _T_2991 | io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 | io_Pctrl_isAdd_C31 | io_Pctrl_isStas_32 |
    io_Pctrl_isStsa_32 ? _T_2999 : io_Pctrl_adderRes_ori[63:0]; // @[PIDU.scala 863:111 864:27]
  wire [63:0] _GEN_575 = _T_2395 | io_Pctrl_isAdd_Q15 | io_Pctrl_isSub_Q15 | io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 ?
    _T_2987 : _GEN_574; // @[PIDU.scala 860:90 861:27]
  wire  _T_3010 = _T_297 & (~io_DecodeIn_ctrl_fuOpType[1] | _T_760); // @[PIDU.scala 871:54]
  wire  _T_3025 = (_T_3010 | _T_1712 & (_T_236 & io_DecodeIn_ctrl_func24 | _T_243 & io_DecodeIn_ctrl_func23)) & _T_25; // @[PIDU.scala 872:126]
  wire  _T_3030 = _T_297 | _T_340; // @[PIDU.scala 873:63]
  wire  _T_3036 = _T_3025 | (io_Pctrl_isRs_32 & (_T_297 | _T_340) | io_Pctrl_isLR_32 & io_DecodeIn_ctrl_fuOpType[4]); // @[PIDU.scala 873:21]
  wire  _T_3040 = _T_3036 | io_Pctrl_isLR_Q31 & io_DecodeIn_ctrl_fuOpType[3]; // @[PIDU.scala 874:21]
  wire  _T_3041 = _T_3040 | io_Pctrl_isRs_XLEN; // @[PIDU.scala 875:21]
  MulAdd_onestage MulAdd17_0 ( // @[PIDU.scala 292:28]
    .io_in_srcs_0(MulAdd17_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd17_0_io_in_srcs_1),
    .io_out_result(MulAdd17_0_io_out_result)
  );
  MulAdd_onestage MulAdd17_1 ( // @[PIDU.scala 293:28]
    .io_in_srcs_0(MulAdd17_1_io_in_srcs_0),
    .io_in_srcs_1(MulAdd17_1_io_in_srcs_1),
    .io_out_result(MulAdd17_1_io_out_result)
  );
  MulAdd_onestage_2 MulAdd33_0 ( // @[PIDU.scala 294:28]
    .io_in_srcs_0(MulAdd33_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd33_0_io_in_srcs_1),
    .io_out_result(MulAdd33_0_io_out_result)
  );
  MulAdd_onestage_3 MulAdd65_0 ( // @[PIDU.scala 295:28]
    .io_in_srcs_0(MulAdd65_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd65_0_io_in_srcs_1),
    .io_out_result(MulAdd65_0_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_0 ( // @[PIDU.scala 296:28]
    .io_in_srcs_0(MulAdd9_0_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_0_io_in_srcs_1),
    .io_out_result(MulAdd9_0_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_1 ( // @[PIDU.scala 297:28]
    .io_in_srcs_0(MulAdd9_1_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_1_io_in_srcs_1),
    .io_out_result(MulAdd9_1_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_2 ( // @[PIDU.scala 298:28]
    .io_in_srcs_0(MulAdd9_2_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_2_io_in_srcs_1),
    .io_out_result(MulAdd9_2_io_out_result)
  );
  MulAdd_onestage_4 MulAdd9_3 ( // @[PIDU.scala 299:28]
    .io_in_srcs_0(MulAdd9_3_io_in_srcs_0),
    .io_in_srcs_1(MulAdd9_3_io_in_srcs_1),
    .io_out_result(MulAdd9_3_io_out_result)
  );
  assign io_Pctrl_isAdd_64 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h2 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h0 &
    io_DecodeIn_ctrl_funct3 == 3'h1; // @[PIDU.scala 154:74]
  assign io_Pctrl_isAdd_32 = _T_3 & (io_DecodeIn_ctrl_fuOpType[6:5] == 2'h0 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h4) &
    io_DecodeIn_ctrl_funct3 == 3'h2; // @[PIDU.scala 155:103]
  assign io_Pctrl_isAdd_16 = _T_14 & io_DecodeIn_ctrl_funct3 == 3'h0; // @[PIDU.scala 156:103]
  assign io_Pctrl_isAdd_8 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h4 & _T_13 & _T_25; // @[PIDU.scala 157:103]
  assign io_Pctrl_isAdd_Q15 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h0 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h2 & _T_5; // @[PIDU.scala 158:75]
  assign io_Pctrl_isAdd_Q31 = _T_38 & _T_3 & _T_5; // @[PIDU.scala 159:75]
  assign io_Pctrl_isAdd_C31 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h1 & _T_3 & _T_5; // @[PIDU.scala 160:75]
  assign io_Pctrl_isAve = io_DecodeIn_ctrl_fuOpType == 7'h70 & _T_25; // @[PIDU.scala 161:48]
  assign io_Pctrl_isAdd = io_Pctrl_isAdd_64 | io_Pctrl_isAdd_32 | io_Pctrl_isAdd_16 | io_Pctrl_isAdd_8 |
    io_Pctrl_isAdd_Q15 | io_Pctrl_isAdd_Q31 | io_Pctrl_isAdd_C31 | io_Pctrl_isAve; // @[PIDU.scala 162:163]
  assign io_Pctrl_isSub_64 = _T_1 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h1 & _T_5; // @[PIDU.scala 164:74]
  assign io_Pctrl_isSub_32 = _T_71 & _T_13 & _T_15; // @[PIDU.scala 165:103]
  assign io_Pctrl_isSub_16 = _T_82 & _T_25; // @[PIDU.scala 166:103]
  assign io_Pctrl_isSub_8 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h5 & _T_13 & _T_25; // @[PIDU.scala 167:103]
  assign io_Pctrl_isSub_Q15 = _T_38 & io_DecodeIn_ctrl_fuOpType[2:0] == 3'h3 & _T_5; // @[PIDU.scala 168:75]
  assign io_Pctrl_isSub_Q31 = _T_38 & _T_71 & _T_5; // @[PIDU.scala 169:75]
  assign io_Pctrl_isSub_C31 = _T_52 & _T_71 & _T_5; // @[PIDU.scala 170:75]
  assign io_Pctrl_isCras_16 = _T_40 & _T_13 & _T_25; // @[PIDU.scala 172:103]
  assign io_Pctrl_isCrsa_16 = _T_108 & _T_13 & _T_25; // @[PIDU.scala 173:103]
  assign io_Pctrl_isCras_32 = _T_133 & _T_15; // @[PIDU.scala 174:103]
  assign io_Pctrl_isCrsa_32 = _T_143 & _T_15; // @[PIDU.scala 175:103]
  assign io_Pctrl_isCr = io_Pctrl_isCras_16 | io_Pctrl_isCrsa_16 | io_Pctrl_isCras_32 | io_Pctrl_isCrsa_32; // @[PIDU.scala 176:83]
  assign io_Pctrl_isStas_16 = (io_DecodeIn_ctrl_fuOpType[6:5] == 2'h3 | io_DecodeIn_ctrl_fuOpType[6:4] == 3'h5) & _T_40
     & _T_15; // @[PIDU.scala 178:103]
  assign io_Pctrl_isStsa_16 = _T_173 & _T_108 & _T_15; // @[PIDU.scala 179:103]
  assign io_Pctrl_isStas_32 = _T_173 & _T_3 & _T_15; // @[PIDU.scala 180:103]
  assign io_Pctrl_isStsa_32 = _T_173 & _T_71 & _T_15; // @[PIDU.scala 181:103]
  assign io_Pctrl_isSt = io_Pctrl_isStas_16 | io_Pctrl_isStsa_16 | io_Pctrl_isStas_32 | io_Pctrl_isStsa_32; // @[PIDU.scala 182:83]
  assign io_Pctrl_isComp_16 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h6 & _T_13 & _T_25; // @[PIDU.scala 184:96]
  assign io_Pctrl_isComp_8 = io_DecodeIn_ctrl_fuOpType[2:0] == 3'h7 & _T_13 & _T_25; // @[PIDU.scala 185:96]
  assign io_Pctrl_isCompare = io_Pctrl_isComp_16 | io_Pctrl_isComp_8; // @[PIDU.scala 186:46]
  assign io_Pctrl_isMaxMin_16 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h4 & io_DecodeIn_ctrl_fuOpType[2:1] == 2'h0 & _T_25; // @[PIDU.scala 188:69]
  assign io_Pctrl_isMaxMin_8 = _T_234 & io_DecodeIn_ctrl_fuOpType[2:1] == 2'h2 & _T_25; // @[PIDU.scala 189:69]
  assign io_Pctrl_isMaxMin_XLEN = io_DecodeIn_ctrl_fuOpType == 7'h5 & io_DecodeIn_ctrl_funct3[2] & ~
    io_DecodeIn_ctrl_funct3[0] & io_DecodeIn_cf_instr[6:0] == 7'h33; // @[PIDU.scala 190:101]
  assign io_Pctrl_isMaxMin_32 = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h9 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'ha) &
    _T_236 & _T_15; // @[PIDU.scala 191:104]
  assign io_Pctrl_isMaxMin = io_Pctrl_isMaxMin_16 | io_Pctrl_isMaxMin_8 | io_Pctrl_isMaxMin_XLEN | io_Pctrl_isMaxMin_32; // @[PIDU.scala 192:98]
  assign io_Pctrl_isPbs = io_DecodeIn_ctrl_fuOpType[6:1] == 6'h3f & _T_25; // @[PIDU.scala 194:53]
  assign io_Pctrl_isRs_16 = io_DecodeIn_ctrl_fuOpType[6:5] == 2'h1 & io_DecodeIn_ctrl_fuOpType[4:3] != 2'h0 & _T_236 &
    _T_25; // @[PIDU.scala 196:85]
  assign io_Pctrl_isLs_16 = _T_278 & _T_40 & _T_25; // @[PIDU.scala 197:85]
  assign io_Pctrl_isLR_16 = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h5 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h6) & _T_108
     & _T_25; // @[PIDU.scala 198:85]
  assign io_Pctrl_isRs_8 = _T_278 & _T_243 & _T_25; // @[PIDU.scala 199:85]
  assign io_Pctrl_isLs_8 = _T_278 & _T_213 & _T_25; // @[PIDU.scala 200:85]
  assign io_Pctrl_isLR_8 = _T_298 & _T_223 & _T_25; // @[PIDU.scala 201:85]
  assign io_Pctrl_isRs_32 = (_T_278 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h8) & _T_236 & _T_15; // @[PIDU.scala 202:111]
  assign io_Pctrl_isLs_32 = _T_341 & _T_40 & _T_15; // @[PIDU.scala 203:111]
  assign io_Pctrl_isLR_32 = _T_301 & _T_15; // @[PIDU.scala 204:86]
  assign io_Pctrl_isLR_Q31 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h3 & _T_223 & _T_5; // @[PIDU.scala 205:74]
  assign io_Pctrl_isLs_Q31 = _T_52 & _T_108 & _T_5; // @[PIDU.scala 206:74]
  assign io_Pctrl_isRs_XLEN = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h2 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'hd) &
    io_DecodeIn_ctrl_fuOpType[2:1] == 2'h1 & _T_5; // @[PIDU.scala 207:103]
  assign io_Pctrl_isSRAIWU = io_DecodeIn_ctrl_fuOpType == 7'h1a & _T_5; // @[PIDU.scala 208:47]
  assign io_Pctrl_isFSRW = io_DecodeIn_cf_instr[26:25] == 2'h2 & io_DecodeIn_ctrl_funct3 == 3'h5 &
    io_DecodeIn_ctrl_fuOpType == 7'h3b; // @[PIDU.scala 209:91]
  assign io_Pctrl_isWext = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h6 & _T_223 & _T_25; // @[PIDU.scala 210:76]
  assign io_Pctrl_isShifter = io_Pctrl_isRs_16 | io_Pctrl_isLs_16 | io_Pctrl_isLR_16 | io_Pctrl_isRs_8 | io_Pctrl_isLs_8
     | io_Pctrl_isLR_8 | io_Pctrl_isRs_32 | io_Pctrl_isLs_32 | io_Pctrl_isLR_32 | io_Pctrl_isLs_Q31 | io_Pctrl_isLR_Q31
     | io_Pctrl_isRs_XLEN | io_Pctrl_isSRAIWU | io_Pctrl_isFSRW | io_Pctrl_isWext; // @[PIDU.scala 211:292]
  assign io_Pctrl_isClip_16 = io_DecodeIn_ctrl_fuOpType == 7'h42 & _T_25; // @[PIDU.scala 213:49]
  assign io_Pctrl_isClip_8 = io_DecodeIn_ctrl_fuOpType == 7'h46 & _T_25; // @[PIDU.scala 214:49]
  assign io_Pctrl_isclip_32 = io_DecodeIn_ctrl_fuOpType[6:4] == 3'h7 & _T_40 & _T_25; // @[PIDU.scala 215:75]
  assign io_Pctrl_isClip = io_Pctrl_isClip_16 | io_Pctrl_isClip_8 | io_Pctrl_isclip_32; // @[PIDU.scala 216:66]
  assign io_Pctrl_isSat_16 = io_DecodeIn_ctrl_fuOpType == 7'h56 & io_DecodeIn_data_src2[4:0] == 5'h11 & _T_25; // @[PIDU.scala 218:77]
  assign io_Pctrl_isSat_8 = _T_439 & io_DecodeIn_data_src2[4:0] == 5'h10 & _T_25; // @[PIDU.scala 219:77]
  assign io_Pctrl_isSat_32 = _T_439 & io_DecodeIn_data_src2[4:0] == 5'h12 & _T_25; // @[PIDU.scala 220:77]
  assign io_Pctrl_isSat_W = _T_439 & io_DecodeIn_data_src2[4:0] == 5'h14 & _T_25; // @[PIDU.scala 221:77]
  assign io_Pctrl_isSat = io_Pctrl_isSat_16 | io_Pctrl_isSat_8 | io_Pctrl_isSat_32 | io_Pctrl_isSat_W; // @[PIDU.scala 222:84]
  assign io_Pctrl_isCnt_16 = io_DecodeIn_ctrl_fuOpType == 7'h57 & io_DecodeIn_data_src2[4:1] == 4'h4 & _T_25; // @[PIDU.scala 224:76]
  assign io_Pctrl_isCnt_8 = _T_466 & io_DecodeIn_data_src2[4:1] == 4'h0 & _T_25; // @[PIDU.scala 225:76]
  assign io_Pctrl_isCnt_32 = _T_466 & io_DecodeIn_data_src2[4:1] == 4'hc & _T_25; // @[PIDU.scala 226:76]
  assign io_Pctrl_isCnt = io_Pctrl_isCnt_16 | io_Pctrl_isCnt_8 | io_Pctrl_isCnt_32; // @[PIDU.scala 227:64]
  assign io_Pctrl_isSwap_16 = _T_10 & _T_223 & _T_5; // @[PIDU.scala 229:72]
  assign io_Pctrl_isSwap_8 = _T_439 & (io_DecodeIn_data_src2[4:0] == 5'h18 & _T_25 & io_DecodeIn_cf_instrType == 5'h15
     | io_DecodeIn_data_src2[5:0] == 6'h8 & _T_399 & io_DecodeIn_cf_instrType == 5'h17); // @[PIDU.scala 230:49]
  assign io_Pctrl_isSwap = io_Pctrl_isSwap_16 | io_Pctrl_isSwap_8; // @[PIDU.scala 231:46]
  assign io_Pctrl_isUnpack = _T_439 & (io_DecodeIn_data_src2[4:3] == 2'h1 | io_DecodeIn_data_src2[4:0] == 5'h13 |
    io_DecodeIn_data_src2[4:0] == 5'h17) & _T_25; // @[PIDU.scala 233:132]
  assign io_Pctrl_isBitrev = _T_530 | io_DecodeIn_ctrl_fuOpType == 7'h35 & _T_399 & io_DecodeIn_cf_instr[6:0] == 7'h13
     & io_DecodeIn_data_src2[4:0] == 5'h1f; // @[PIDU.scala 236:24]
  assign io_Pctrl_isCmix = io_DecodeIn_cf_instr[14:12] == 3'h1 & _T_255 & io_DecodeIn_cf_instr[26:25] == 2'h3; // @[PIDU.scala 238:114]
  assign io_Pctrl_isInsertb = _T_439 & io_DecodeIn_cf_instr[24:23] == 2'h0 & _T_25; // @[PIDU.scala 240:92]
  assign io_Pctrl_isPackbb = io_DecodeIn_ctrl_fuOpType == 7'h4 & io_DecodeIn_ctrl_funct3 == 3'h4 & _T_255; // @[PIDU.scala 242:72]
  assign io_Pctrl_isPackbt = io_DecodeIn_ctrl_fuOpType == 7'hf & _T_15; // @[PIDU.scala 243:49]
  assign io_Pctrl_isPacktb = io_DecodeIn_ctrl_fuOpType == 7'h1f & _T_15; // @[PIDU.scala 244:49]
  assign io_Pctrl_isPacktt = io_DecodeIn_ctrl_fuOpType == 7'h24 & _T_556 & _T_255; // @[PIDU.scala 245:72]
  assign io_Pctrl_isPack = io_Pctrl_isPackbb | io_Pctrl_isPackbt | io_Pctrl_isPacktb | io_Pctrl_isPacktt; // @[PIDU.scala 246:85]
  assign io_Pctrl_isSub = _T_1748 | io_Pctrl_isComp_8 | io_Pctrl_isMaxMin | io_Pctrl_isPbs | io_Pctrl_isSub_Q15 |
    io_Pctrl_isSub_Q31 | io_Pctrl_isSub_C31 ? 8'hff : {{4'd0}, _GEN_379}; // @[PIDU.scala 634:125 635:23]
  assign io_Pctrl_isAdder = (io_Pctrl_isSub != 8'h0 | io_Pctrl_isAdd | io_Pctrl_isCr | io_Pctrl_isSt) & ~
    io_Pctrl_isCompare & ~io_Pctrl_isMaxMin & ~io_Pctrl_isPbs; // @[PIDU.scala 646:142]
  assign io_Pctrl_SrcSigned = _T_38 | _T_234 | io_Pctrl_isSt & (io_DecodeIn_ctrl_fuOpType[6:3] == 4'hb | _T_633); // @[PIDU.scala 648:73]
  assign io_Pctrl_Saturating = ~io_Pctrl_isSt & io_DecodeIn_ctrl_fuOpType[3] | io_Pctrl_isSt & ~
    io_DecodeIn_ctrl_fuOpType[3]; // @[PIDU.scala 649:62]
  assign io_Pctrl_Translation = ~io_Pctrl_Saturating & (_T_1781 & ~_T_12 | io_Pctrl_isSt & (_T_1775 | _T_387)); // @[PIDU.scala 650:50]
  assign io_Pctrl_LessEqual = io_Pctrl_Saturating; // @[PIDU.scala 651:26]
  assign io_Pctrl_LessThan = io_Pctrl_Translation; // @[PIDU.scala 652:26]
  assign io_Pctrl_adderRes_ori = _T_2955[79:0]; // @[PIDU.scala 840:27]
  assign io_Pctrl_adderRes = _T_1804 | io_Pctrl_isPbs ? _T_2973 : _GEN_575; // @[PIDU.scala 857:65 858:27]
  assign io_Pctrl_adderRes_ori_drophighestbit = _T_2956[79:0]; // @[PIDU.scala 841:42]
  assign io_Pctrl_Round = _T_3041 | io_Pctrl_isSRAIWU; // @[PIDU.scala 876:21]
  assign io_Pctrl_ShiftSigned = io_Pctrl_isLR_16 | io_Pctrl_isLR_8 | io_Pctrl_isLR_32 | io_Pctrl_isLR_Q31 |
    io_Pctrl_isLs_Q31 | io_Pctrl_isLs_32 & _T_3030 | (io_Pctrl_isLs_16 | io_Pctrl_isLs_8) & (_T_297 |
    io_DecodeIn_ctrl_fuOpType == 7'h3a & io_DecodeIn_ctrl_func24 | _T_1288 & io_DecodeIn_ctrl_func23); // @[PIDU.scala 877:191]
  assign io_Pctrl_Arithmetic = (io_Pctrl_isRs_16 | io_Pctrl_isRs_8 | io_Pctrl_isRs_32) & ~io_DecodeIn_ctrl_fuOpType[0]
     | io_Pctrl_isLR_16 | io_Pctrl_isLR_8 | io_Pctrl_isLR_32 | io_Pctrl_isLR_Q31 | io_Pctrl_isRs_XLEN |
    io_Pctrl_isSRAIWU; // @[PIDU.scala 878:209]
  assign io_Pctrl_isMul_16 = ~io_DecodeIn_ctrl_fuOpType[2] & _T_25; // @[PIDU.scala 248:43]
  assign io_Pctrl_isMul_8 = io_DecodeIn_ctrl_fuOpType[2] & _T_25 & io_DecodeIn_ctrl_fuOpType[6:3] != 4'hc; // @[PIDU.scala 249:61]
  assign io_Pctrl_isMSW_3232 = _T_275 & _T_236 & _T_5; // @[PIDU.scala 250:76]
  assign io_Pctrl_isMSW_3216 = (_T_275 & _T_390 | io_DecodeIn_ctrl_fuOpType[6] & _T_223) & _T_5; // @[PIDU.scala 251:126]
  assign io_Pctrl_isS1632 = ~io_DecodeIn_ctrl_fuOpType[6] & (_T_28 | _T_96 & io_DecodeIn_ctrl_fuOpType[6:3] > 4'h2 |
    _T_213 & io_DecodeIn_ctrl_fuOpType[5] | io_DecodeIn_ctrl_fuOpType == 7'h27) & _T_5; // @[PIDU.scala 252:187]
  assign io_Pctrl_isS1664 = io_DecodeIn_ctrl_fuOpType == 7'h2f & _T_5; // @[PIDU.scala 253:49]
  assign io_Pctrl_is832 = io_DecodeIn_ctrl_fuOpType[6:3] == 4'hc & io_DecodeIn_ctrl_fuOpType[2:0] != 3'h7 & _T_25; // @[PIDU.scala 254:77]
  assign io_Pctrl_is3264 = _T_1 & _T_390 & _T_5; // @[PIDU.scala 255:74]
  assign io_Pctrl_is1664 = _T_1 & _T_635 & _T_5; // @[PIDU.scala 256:75]
  assign io_Pctrl_isQ15orQ31 = (_T_10 & (_T_213 | _T_96) | _T_170 & _T_71 & _T_277) & _T_5; // @[PIDU.scala 257:183]
  assign io_Pctrl_isC31 = (_T_431 & _T_3 | _T_633 & _T_390) & _T_5; // @[PIDU.scala 258:130]
  assign io_Pctrl_isQ15_64ONLY = _T_170 & _T_277 & io_DecodeIn_ctrl_fuOpType[2] & io_DecodeIn_ctrl_fuOpType[1:0] != 2'h3
     & _T_5; // @[PIDU.scala 259:123]
  assign io_Pctrl_isQ63_64ONLY = _T_278 & _T_96 & _T_15; // @[PIDU.scala 260:102]
  assign io_Pctrl_isMul_32_64ONLY = (_T_385 | io_DecodeIn_ctrl_fuOpType[6:3] == 4'h1) & _T_28 & _T_15; // @[PIDU.scala 261:113]
  assign io_Pctrl_isPMA_64ONLY = (io_DecodeIn_ctrl_fuOpType[6:3] == 4'h3 & _T_243 | _T_12 & io_DecodeIn_ctrl_fuOpType[2]
     | (_T_28 | _T_213) & _T_275 & _T_277) & _T_15; // @[PIDU.scala 262:223]
  assign io_Pctrl_mulres9_0 = MulAdd9_0_io_out_result; // @[PIDU.scala 622:25]
  assign io_Pctrl_mulres9_1 = MulAdd9_1_io_out_result; // @[PIDU.scala 623:25]
  assign io_Pctrl_mulres9_2 = MulAdd9_2_io_out_result; // @[PIDU.scala 624:25]
  assign io_Pctrl_mulres9_3 = MulAdd9_3_io_out_result; // @[PIDU.scala 625:25]
  assign io_Pctrl_mulres17_0 = MulAdd17_0_io_out_result; // @[PIDU.scala 626:25]
  assign io_Pctrl_mulres17_1 = MulAdd17_1_io_out_result; // @[PIDU.scala 627:25]
  assign io_Pctrl_mulres33_0 = MulAdd33_0_io_out_result; // @[PIDU.scala 628:25]
  assign io_Pctrl_mulres65_0 = MulAdd65_0_io_out_result; // @[PIDU.scala 629:25]
  assign MulAdd17_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? _GEN_22 : _GEN_332; // @[PIDU.scala 311:32]
  assign MulAdd17_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? _GEN_26 : _GEN_340; // @[PIDU.scala 311:32]
  assign MulAdd17_1_io_in_srcs_0 = _GEN_353[16:0];
  assign MulAdd17_1_io_in_srcs_1 = _GEN_357[16:0];
  assign MulAdd33_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? _GEN_24 : _GEN_334; // @[PIDU.scala 311:32]
  assign MulAdd33_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? _GEN_28 : _GEN_342; // @[PIDU.scala 311:32]
  assign MulAdd65_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? _GEN_25 : _GEN_335; // @[PIDU.scala 311:32]
  assign MulAdd65_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? _GEN_29 : _GEN_343; // @[PIDU.scala 311:32]
  assign MulAdd9_0_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_328; // @[PIDU.scala 305:22 311:32]
  assign MulAdd9_0_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_336; // @[PIDU.scala 305:22 311:32]
  assign MulAdd9_1_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_329; // @[PIDU.scala 306:22 311:32]
  assign MulAdd9_1_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_337; // @[PIDU.scala 306:22 311:32]
  assign MulAdd9_2_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_330; // @[PIDU.scala 307:22 311:32]
  assign MulAdd9_2_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_338; // @[PIDU.scala 307:22 311:32]
  assign MulAdd9_3_io_in_srcs_0 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_331; // @[PIDU.scala 308:22 311:32]
  assign MulAdd9_3_io_in_srcs_1 = io_Pctrl_isMul_16 ? 9'h0 : _GEN_339; // @[PIDU.scala 308:22 311:32]
endmodule
module SIMDU_2way(
  input         clock,
  input         reset,
  input         io_flush,
  output [38:0] io_DecodeOut_0_cf_pc,
  output [63:0] io_DecodeOut_0_cf_runahead_checkpoint_id,
  output        io_DecodeOut_0_ctrl_rfWen,
  output [4:0]  io_DecodeOut_0_ctrl_rfDest,
  output        io_DecodeOut_0_pext_OV,
  output [4:0]  io_DecodeOut_0_InstNo,
  output [38:0] io_DecodeOut_1_cf_pc,
  output [63:0] io_DecodeOut_1_cf_runahead_checkpoint_id,
  output        io_DecodeOut_1_ctrl_rfWen,
  output [4:0]  io_DecodeOut_1_ctrl_rfDest,
  output        io_DecodeOut_1_pext_OV,
  output [4:0]  io_DecodeOut_1_InstNo,
  input  [63:0] io_DecodeIn_0_cf_instr,
  input  [38:0] io_DecodeIn_0_cf_pc,
  input  [63:0] io_DecodeIn_0_cf_runahead_checkpoint_id,
  input  [4:0]  io_DecodeIn_0_cf_instrType,
  input  [6:0]  io_DecodeIn_0_ctrl_fuOpType,
  input  [2:0]  io_DecodeIn_0_ctrl_funct3,
  input         io_DecodeIn_0_ctrl_func24,
  input         io_DecodeIn_0_ctrl_func23,
  input         io_DecodeIn_0_ctrl_rfWen,
  input  [4:0]  io_DecodeIn_0_ctrl_rfDest,
  input  [63:0] io_DecodeIn_0_data_src1,
  input  [63:0] io_DecodeIn_0_data_src2,
  input  [63:0] io_DecodeIn_0_data_src3,
  input  [4:0]  io_DecodeIn_0_InstNo,
  input         io_DecodeIn_0_InstFlag,
  input  [63:0] io_DecodeIn_1_cf_instr,
  input  [38:0] io_DecodeIn_1_cf_pc,
  input  [63:0] io_DecodeIn_1_cf_runahead_checkpoint_id,
  input  [4:0]  io_DecodeIn_1_cf_instrType,
  input  [6:0]  io_DecodeIn_1_ctrl_fuOpType,
  input  [2:0]  io_DecodeIn_1_ctrl_funct3,
  input         io_DecodeIn_1_ctrl_func24,
  input         io_DecodeIn_1_ctrl_func23,
  input         io_DecodeIn_1_ctrl_rfWen,
  input  [4:0]  io_DecodeIn_1_ctrl_rfDest,
  input  [63:0] io_DecodeIn_1_data_src1,
  input  [63:0] io_DecodeIn_1_data_src2,
  input  [63:0] io_DecodeIn_1_data_src3,
  input  [4:0]  io_DecodeIn_1_InstNo,
  input         io_DecodeIn_1_InstFlag,
  output        io_FirstStageFire_0,
  output        io_FirstStageFire_1,
  output        io_in_0_ready,
  input         io_in_0_valid,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [63:0] io_out_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [95:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [95:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [95:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [95:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [95:0] _RAND_229;
  reg [159:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [95:0] _RAND_263;
  reg [159:0] _RAND_264;
  reg [31:0] _RAND_265;
`endif // RANDOMIZE_REG_INIT
  wire  PALU0_io_in_ready; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_valid; // @[SIMDU.scala 451:21]
  wire [38:0] PALU0_io_in_bits_DecodeIn_cf_pc; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 451:21]
  wire [6:0] PALU0_io_in_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 451:21]
  wire [2:0] PALU0_io_in_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 451:21]
  wire [4:0] PALU0_io_in_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_in_bits_DecodeIn_data_src1; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_in_bits_DecodeIn_data_src2; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_in_bits_DecodeIn_data_src3; // @[SIMDU.scala 451:21]
  wire [4:0] PALU0_io_in_bits_DecodeIn_InstNo; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_DecodeIn_InstFlag; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_64; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAve; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_64; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSub_C31; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCras_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCras_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isStas_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isStsa_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isStas_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isStsa_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isComp_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isComp_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCompare; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isMaxMin; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isPbs; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isRs_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLs_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLR_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isRs_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLs_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLR_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isRs_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLs_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLR_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isFSRW; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isWext; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isShifter; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isClip_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isClip_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isclip_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isClip; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSat_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSat_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSat_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSat_W; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSat; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCnt_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCnt_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCnt_32; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCnt; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSwap_16; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSwap_8; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isSwap; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isUnpack; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isBitrev; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isCmix; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isInsertb; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isPackbb; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isPackbt; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isPacktb; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isPacktt; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isPack; // @[SIMDU.scala 451:21]
  wire [7:0] PALU0_io_in_bits_Pctrl_isSub; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_isAdder; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_SrcSigned; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_Saturating; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_Translation; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_LessEqual; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_LessThan; // @[SIMDU.scala 451:21]
  wire [79:0] PALU0_io_in_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_in_bits_Pctrl_adderRes; // @[SIMDU.scala 451:21]
  wire [79:0] PALU0_io_in_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_Round; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 451:21]
  wire  PALU0_io_in_bits_Pctrl_Arithmetic; // @[SIMDU.scala 451:21]
  wire  PALU0_io_out_ready; // @[SIMDU.scala 451:21]
  wire  PALU0_io_out_valid; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_out_bits_result; // @[SIMDU.scala 451:21]
  wire [38:0] PALU0_io_out_bits_DecodeOut_cf_pc; // @[SIMDU.scala 451:21]
  wire [63:0] PALU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id; // @[SIMDU.scala 451:21]
  wire  PALU0_io_out_bits_DecodeOut_ctrl_rfWen; // @[SIMDU.scala 451:21]
  wire [4:0] PALU0_io_out_bits_DecodeOut_ctrl_rfDest; // @[SIMDU.scala 451:21]
  wire  PALU0_io_out_bits_DecodeOut_pext_OV; // @[SIMDU.scala 451:21]
  wire [4:0] PALU0_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 451:21]
  wire  PALU0_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 451:21]
  wire  PMDU0_io_in_ready; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_valid; // @[SIMDU.scala 452:21]
  wire [38:0] PMDU0_io_in_bits_DecodeIn_cf_pc; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 452:21]
  wire [6:0] PMDU0_io_in_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 452:21]
  wire [4:0] PMDU0_io_in_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_in_bits_DecodeIn_data_src1; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_in_bits_DecodeIn_data_src2; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_in_bits_DecodeIn_data_src3; // @[SIMDU.scala 452:21]
  wire [4:0] PMDU0_io_in_bits_DecodeIn_InstNo; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_DecodeIn_InstFlag; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isMul_16; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isMul_8; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isS1632; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isS1664; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_is832; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_is3264; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_is1664; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isC31; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_in_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 452:21]
  wire [17:0] PMDU0_io_in_bits_Pctrl_mulres9_0; // @[SIMDU.scala 452:21]
  wire [17:0] PMDU0_io_in_bits_Pctrl_mulres9_1; // @[SIMDU.scala 452:21]
  wire [17:0] PMDU0_io_in_bits_Pctrl_mulres9_2; // @[SIMDU.scala 452:21]
  wire [17:0] PMDU0_io_in_bits_Pctrl_mulres9_3; // @[SIMDU.scala 452:21]
  wire [33:0] PMDU0_io_in_bits_Pctrl_mulres17_0; // @[SIMDU.scala 452:21]
  wire [33:0] PMDU0_io_in_bits_Pctrl_mulres17_1; // @[SIMDU.scala 452:21]
  wire [65:0] PMDU0_io_in_bits_Pctrl_mulres33_0; // @[SIMDU.scala 452:21]
  wire [129:0] PMDU0_io_in_bits_Pctrl_mulres65_0; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_out_ready; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_out_valid; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_out_bits_result; // @[SIMDU.scala 452:21]
  wire [38:0] PMDU0_io_out_bits_DecodeOut_cf_pc; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id; // @[SIMDU.scala 452:21]
  wire [6:0] PMDU0_io_out_bits_DecodeOut_ctrl_fuOpType; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_out_bits_DecodeOut_ctrl_rfWen; // @[SIMDU.scala 452:21]
  wire [4:0] PMDU0_io_out_bits_DecodeOut_ctrl_rfDest; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_out_bits_DecodeOut_data_src1; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_out_bits_DecodeOut_data_src2; // @[SIMDU.scala 452:21]
  wire [63:0] PMDU0_io_out_bits_DecodeOut_data_src3; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_out_bits_DecodeOut_pext_OV; // @[SIMDU.scala 452:21]
  wire [4:0] PMDU0_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 452:21]
  wire  PMDU0_io_FirstStageFire; // @[SIMDU.scala 452:21]
  wire  PALU1_io_in_ready; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_valid; // @[SIMDU.scala 453:21]
  wire [38:0] PALU1_io_in_bits_DecodeIn_cf_pc; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 453:21]
  wire [6:0] PALU1_io_in_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 453:21]
  wire [2:0] PALU1_io_in_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 453:21]
  wire [4:0] PALU1_io_in_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_in_bits_DecodeIn_data_src1; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_in_bits_DecodeIn_data_src2; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_in_bits_DecodeIn_data_src3; // @[SIMDU.scala 453:21]
  wire [4:0] PALU1_io_in_bits_DecodeIn_InstNo; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_DecodeIn_InstFlag; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_64; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAve; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_64; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSub_C31; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCras_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCras_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isStas_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isStsa_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isStas_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isStsa_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isComp_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isComp_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCompare; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isMaxMin; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isPbs; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isRs_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLs_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLR_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isRs_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLs_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLR_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isRs_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLs_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLR_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isFSRW; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isWext; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isShifter; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isClip_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isClip_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isclip_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isClip; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSat_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSat_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSat_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSat_W; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSat; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCnt_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCnt_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCnt_32; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCnt; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSwap_16; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSwap_8; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isSwap; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isUnpack; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isBitrev; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isCmix; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isInsertb; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isPackbb; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isPackbt; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isPacktb; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isPacktt; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isPack; // @[SIMDU.scala 453:21]
  wire [7:0] PALU1_io_in_bits_Pctrl_isSub; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_isAdder; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_SrcSigned; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_Saturating; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_Translation; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_LessEqual; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_LessThan; // @[SIMDU.scala 453:21]
  wire [79:0] PALU1_io_in_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_in_bits_Pctrl_adderRes; // @[SIMDU.scala 453:21]
  wire [79:0] PALU1_io_in_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_Round; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 453:21]
  wire  PALU1_io_in_bits_Pctrl_Arithmetic; // @[SIMDU.scala 453:21]
  wire  PALU1_io_out_ready; // @[SIMDU.scala 453:21]
  wire  PALU1_io_out_valid; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_out_bits_result; // @[SIMDU.scala 453:21]
  wire [38:0] PALU1_io_out_bits_DecodeOut_cf_pc; // @[SIMDU.scala 453:21]
  wire [63:0] PALU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id; // @[SIMDU.scala 453:21]
  wire  PALU1_io_out_bits_DecodeOut_ctrl_rfWen; // @[SIMDU.scala 453:21]
  wire [4:0] PALU1_io_out_bits_DecodeOut_ctrl_rfDest; // @[SIMDU.scala 453:21]
  wire  PALU1_io_out_bits_DecodeOut_pext_OV; // @[SIMDU.scala 453:21]
  wire [4:0] PALU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 453:21]
  wire  PALU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 453:21]
  wire  PMDU1_io_in_ready; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_valid; // @[SIMDU.scala 454:21]
  wire [38:0] PMDU1_io_in_bits_DecodeIn_cf_pc; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_in_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 454:21]
  wire [6:0] PMDU1_io_in_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 454:21]
  wire [4:0] PMDU1_io_in_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_in_bits_DecodeIn_data_src1; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_in_bits_DecodeIn_data_src2; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_in_bits_DecodeIn_data_src3; // @[SIMDU.scala 454:21]
  wire [4:0] PMDU1_io_in_bits_DecodeIn_InstNo; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_DecodeIn_InstFlag; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isMul_16; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isMul_8; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isS1632; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isS1664; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_is832; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_is3264; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_is1664; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isC31; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_in_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 454:21]
  wire [17:0] PMDU1_io_in_bits_Pctrl_mulres9_0; // @[SIMDU.scala 454:21]
  wire [17:0] PMDU1_io_in_bits_Pctrl_mulres9_1; // @[SIMDU.scala 454:21]
  wire [17:0] PMDU1_io_in_bits_Pctrl_mulres9_2; // @[SIMDU.scala 454:21]
  wire [17:0] PMDU1_io_in_bits_Pctrl_mulres9_3; // @[SIMDU.scala 454:21]
  wire [33:0] PMDU1_io_in_bits_Pctrl_mulres17_0; // @[SIMDU.scala 454:21]
  wire [33:0] PMDU1_io_in_bits_Pctrl_mulres17_1; // @[SIMDU.scala 454:21]
  wire [65:0] PMDU1_io_in_bits_Pctrl_mulres33_0; // @[SIMDU.scala 454:21]
  wire [129:0] PMDU1_io_in_bits_Pctrl_mulres65_0; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_out_ready; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_out_valid; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_out_bits_result; // @[SIMDU.scala 454:21]
  wire [38:0] PMDU1_io_out_bits_DecodeOut_cf_pc; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id; // @[SIMDU.scala 454:21]
  wire [6:0] PMDU1_io_out_bits_DecodeOut_ctrl_fuOpType; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_out_bits_DecodeOut_ctrl_rfWen; // @[SIMDU.scala 454:21]
  wire [4:0] PMDU1_io_out_bits_DecodeOut_ctrl_rfDest; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_out_bits_DecodeOut_data_src1; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_out_bits_DecodeOut_data_src2; // @[SIMDU.scala 454:21]
  wire [63:0] PMDU1_io_out_bits_DecodeOut_data_src3; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_out_bits_DecodeOut_pext_OV; // @[SIMDU.scala 454:21]
  wire [4:0] PMDU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 454:21]
  wire  PMDU1_io_FirstStageFire; // @[SIMDU.scala 454:21]
  wire [63:0] PIDU0_io_DecodeIn_cf_instr; // @[SIMDU.scala 455:21]
  wire [4:0] PIDU0_io_DecodeIn_cf_instrType; // @[SIMDU.scala 455:21]
  wire [6:0] PIDU0_io_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 455:21]
  wire [2:0] PIDU0_io_DecodeIn_ctrl_funct3; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_DecodeIn_ctrl_func24; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_DecodeIn_ctrl_func23; // @[SIMDU.scala 455:21]
  wire [63:0] PIDU0_io_DecodeIn_data_src1; // @[SIMDU.scala 455:21]
  wire [63:0] PIDU0_io_DecodeIn_data_src2; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_64; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_Q15; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_Q31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd_C31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAve; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdd; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_64; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_Q15; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_Q31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSub_C31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCras_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCrsa_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCras_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCrsa_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCr; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isStas_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isStsa_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isStas_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isStsa_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSt; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isComp_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isComp_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCompare; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMaxMin_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMaxMin_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMaxMin_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMaxMin; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPbs; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isRs_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLs_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLR_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isRs_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLs_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLR_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isRs_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLs_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLR_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLR_Q31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isLs_Q31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isRs_XLEN; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSRAIWU; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isFSRW; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isWext; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isShifter; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isClip_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isClip_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isclip_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isClip; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSat_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSat_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSat_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSat_W; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSat; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCnt_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCnt_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCnt_32; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCnt; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSwap_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSwap_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isSwap; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isUnpack; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isBitrev; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isCmix; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isInsertb; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPackbb; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPackbt; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPacktb; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPacktt; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPack; // @[SIMDU.scala 455:21]
  wire [7:0] PIDU0_io_Pctrl_isSub; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isAdder; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_SrcSigned; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_Saturating; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_Translation; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_LessEqual; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_LessThan; // @[SIMDU.scala 455:21]
  wire [79:0] PIDU0_io_Pctrl_adderRes_ori; // @[SIMDU.scala 455:21]
  wire [63:0] PIDU0_io_Pctrl_adderRes; // @[SIMDU.scala 455:21]
  wire [79:0] PIDU0_io_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_Round; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_ShiftSigned; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_Arithmetic; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMul_16; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMul_8; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMSW_3232; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMSW_3216; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isS1632; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isS1664; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_is832; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_is3264; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_is1664; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isQ15orQ31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isC31; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 455:21]
  wire  PIDU0_io_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 455:21]
  wire [17:0] PIDU0_io_Pctrl_mulres9_0; // @[SIMDU.scala 455:21]
  wire [17:0] PIDU0_io_Pctrl_mulres9_1; // @[SIMDU.scala 455:21]
  wire [17:0] PIDU0_io_Pctrl_mulres9_2; // @[SIMDU.scala 455:21]
  wire [17:0] PIDU0_io_Pctrl_mulres9_3; // @[SIMDU.scala 455:21]
  wire [33:0] PIDU0_io_Pctrl_mulres17_0; // @[SIMDU.scala 455:21]
  wire [33:0] PIDU0_io_Pctrl_mulres17_1; // @[SIMDU.scala 455:21]
  wire [65:0] PIDU0_io_Pctrl_mulres33_0; // @[SIMDU.scala 455:21]
  wire [129:0] PIDU0_io_Pctrl_mulres65_0; // @[SIMDU.scala 455:21]
  wire [63:0] PIDU1_io_DecodeIn_cf_instr; // @[SIMDU.scala 456:21]
  wire [4:0] PIDU1_io_DecodeIn_cf_instrType; // @[SIMDU.scala 456:21]
  wire [6:0] PIDU1_io_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 456:21]
  wire [2:0] PIDU1_io_DecodeIn_ctrl_funct3; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_DecodeIn_ctrl_func24; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_DecodeIn_ctrl_func23; // @[SIMDU.scala 456:21]
  wire [63:0] PIDU1_io_DecodeIn_data_src1; // @[SIMDU.scala 456:21]
  wire [63:0] PIDU1_io_DecodeIn_data_src2; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_64; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_Q15; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_Q31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd_C31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAve; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdd; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_64; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_Q15; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_Q31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSub_C31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCras_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCrsa_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCras_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCrsa_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCr; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isStas_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isStsa_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isStas_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isStsa_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSt; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isComp_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isComp_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCompare; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMaxMin_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMaxMin_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMaxMin_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMaxMin; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPbs; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isRs_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLs_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLR_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isRs_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLs_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLR_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isRs_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLs_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLR_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLR_Q31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isLs_Q31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isRs_XLEN; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSRAIWU; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isFSRW; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isWext; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isShifter; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isClip_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isClip_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isclip_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isClip; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSat_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSat_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSat_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSat_W; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSat; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCnt_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCnt_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCnt_32; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCnt; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSwap_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSwap_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isSwap; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isUnpack; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isBitrev; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isCmix; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isInsertb; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPackbb; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPackbt; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPacktb; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPacktt; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPack; // @[SIMDU.scala 456:21]
  wire [7:0] PIDU1_io_Pctrl_isSub; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isAdder; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_SrcSigned; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_Saturating; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_Translation; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_LessEqual; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_LessThan; // @[SIMDU.scala 456:21]
  wire [79:0] PIDU1_io_Pctrl_adderRes_ori; // @[SIMDU.scala 456:21]
  wire [63:0] PIDU1_io_Pctrl_adderRes; // @[SIMDU.scala 456:21]
  wire [79:0] PIDU1_io_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_Round; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_ShiftSigned; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_Arithmetic; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMul_16; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMul_8; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMSW_3232; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMSW_3216; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isS1632; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isS1664; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_is832; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_is3264; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_is1664; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isQ15orQ31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isC31; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 456:21]
  wire  PIDU1_io_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 456:21]
  wire [17:0] PIDU1_io_Pctrl_mulres9_0; // @[SIMDU.scala 456:21]
  wire [17:0] PIDU1_io_Pctrl_mulres9_1; // @[SIMDU.scala 456:21]
  wire [17:0] PIDU1_io_Pctrl_mulres9_2; // @[SIMDU.scala 456:21]
  wire [17:0] PIDU1_io_Pctrl_mulres9_3; // @[SIMDU.scala 456:21]
  wire [33:0] PIDU1_io_Pctrl_mulres17_0; // @[SIMDU.scala 456:21]
  wire [33:0] PIDU1_io_Pctrl_mulres17_1; // @[SIMDU.scala 456:21]
  wire [65:0] PIDU1_io_Pctrl_mulres33_0; // @[SIMDU.scala 456:21]
  wire [129:0] PIDU1_io_Pctrl_mulres65_0; // @[SIMDU.scala 456:21]
  reg [38:0] PALU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 482:32]
  reg [63:0] PALU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 482:32]
  reg [6:0] PALU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 482:32]
  reg [2:0] PALU0_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 482:32]
  reg [4:0] PALU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 482:32]
  reg [63:0] PALU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 482:32]
  reg [63:0] PALU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 482:32]
  reg [63:0] PALU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 482:32]
  reg [4:0] PALU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_64; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAve; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_64; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSub_C31; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCras_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCras_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isStas_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isStsa_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isStas_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isStsa_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isComp_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isComp_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCompare; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isMaxMin; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isPbs; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isRs_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLs_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLR_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isRs_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLs_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLR_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isRs_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLs_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLR_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isFSRW; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isWext; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isShifter; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isClip_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isClip_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isclip_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isClip; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSat_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSat_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSat_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSat_W; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSat; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCnt_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCnt_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCnt_32; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCnt; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSwap_16; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSwap_8; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isSwap; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isUnpack; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isBitrev; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isCmix; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isInsertb; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isPackbb; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isPackbt; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isPacktb; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isPacktt; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isPack; // @[SIMDU.scala 482:32]
  reg [7:0] PALU0_bits_Pctrl_isSub; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_isAdder; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_SrcSigned; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_Saturating; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_Translation; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_LessEqual; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_LessThan; // @[SIMDU.scala 482:32]
  reg [79:0] PALU0_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 482:32]
  reg [63:0] PALU0_bits_Pctrl_adderRes; // @[SIMDU.scala 482:32]
  reg [79:0] PALU0_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_Round; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 482:32]
  reg  PALU0_bits_Pctrl_Arithmetic; // @[SIMDU.scala 482:32]
  reg  PALU0_valid; // @[SIMDU.scala 484:28]
  wire  _T_4 = PALU0_io_out_ready & PALU0_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T_4 ? 1'h0 : PALU0_valid; // @[SIMDU.scala 486:19 487:{28,46}]
  reg [38:0] PALU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 490:32]
  reg [63:0] PALU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 490:32]
  reg [6:0] PALU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 490:32]
  reg [2:0] PALU1_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 490:32]
  reg [4:0] PALU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 490:32]
  reg [63:0] PALU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 490:32]
  reg [63:0] PALU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 490:32]
  reg [63:0] PALU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 490:32]
  reg [4:0] PALU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_64; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAve; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_64; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSub_C31; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCras_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCras_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isStas_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isStsa_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isStas_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isStsa_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isComp_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isComp_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCompare; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isMaxMin; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isPbs; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isRs_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLs_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLR_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isRs_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLs_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLR_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isRs_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLs_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLR_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isFSRW; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isWext; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isShifter; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isClip_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isClip_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isclip_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isClip; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSat_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSat_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSat_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSat_W; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSat; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCnt_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCnt_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCnt_32; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCnt; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSwap_16; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSwap_8; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isSwap; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isUnpack; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isBitrev; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isCmix; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isInsertb; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isPackbb; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isPackbt; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isPacktb; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isPacktt; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isPack; // @[SIMDU.scala 490:32]
  reg [7:0] PALU1_bits_Pctrl_isSub; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_isAdder; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_SrcSigned; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_Saturating; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_Translation; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_LessEqual; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_LessThan; // @[SIMDU.scala 490:32]
  reg [79:0] PALU1_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 490:32]
  reg [63:0] PALU1_bits_Pctrl_adderRes; // @[SIMDU.scala 490:32]
  reg [79:0] PALU1_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_Round; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 490:32]
  reg  PALU1_bits_Pctrl_Arithmetic; // @[SIMDU.scala 490:32]
  reg  PALU1_valid; // @[SIMDU.scala 492:28]
  wire  _T_5 = PALU1_io_out_ready & PALU1_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_5 ? 1'h0 : PALU1_valid; // @[SIMDU.scala 494:19 495:{28,46}]
  reg [38:0] PMDU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 499:32]
  reg [63:0] PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 499:32]
  reg [6:0] PMDU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 499:32]
  reg [4:0] PMDU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 499:32]
  reg [63:0] PMDU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 499:32]
  reg [63:0] PMDU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 499:32]
  reg [63:0] PMDU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 499:32]
  reg [4:0] PMDU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isMul_16; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isMul_8; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isS1632; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isS1664; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_is832; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_is3264; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_is1664; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isC31; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 499:32]
  reg  PMDU0_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 499:32]
  reg [17:0] PMDU0_bits_Pctrl_mulres9_0; // @[SIMDU.scala 499:32]
  reg [17:0] PMDU0_bits_Pctrl_mulres9_1; // @[SIMDU.scala 499:32]
  reg [17:0] PMDU0_bits_Pctrl_mulres9_2; // @[SIMDU.scala 499:32]
  reg [17:0] PMDU0_bits_Pctrl_mulres9_3; // @[SIMDU.scala 499:32]
  reg [33:0] PMDU0_bits_Pctrl_mulres17_0; // @[SIMDU.scala 499:32]
  reg [33:0] PMDU0_bits_Pctrl_mulres17_1; // @[SIMDU.scala 499:32]
  reg [65:0] PMDU0_bits_Pctrl_mulres33_0; // @[SIMDU.scala 499:32]
  reg [129:0] PMDU0_bits_Pctrl_mulres65_0; // @[SIMDU.scala 499:32]
  reg  PMDU0_valid; // @[SIMDU.scala 501:28]
  wire  _GEN_2 = PMDU0_io_FirstStageFire ? 1'h0 : PMDU0_valid; // @[SIMDU.scala 503:19 504:{32,50}]
  reg [38:0] PMDU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 507:32]
  reg [63:0] PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 507:32]
  reg [6:0] PMDU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 507:32]
  reg [4:0] PMDU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 507:32]
  reg [63:0] PMDU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 507:32]
  reg [63:0] PMDU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 507:32]
  reg [63:0] PMDU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 507:32]
  reg [4:0] PMDU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isMul_16; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isMul_8; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isS1632; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isS1664; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_is832; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_is3264; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_is1664; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isC31; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 507:32]
  reg  PMDU1_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 507:32]
  reg [17:0] PMDU1_bits_Pctrl_mulres9_0; // @[SIMDU.scala 507:32]
  reg [17:0] PMDU1_bits_Pctrl_mulres9_1; // @[SIMDU.scala 507:32]
  reg [17:0] PMDU1_bits_Pctrl_mulres9_2; // @[SIMDU.scala 507:32]
  reg [17:0] PMDU1_bits_Pctrl_mulres9_3; // @[SIMDU.scala 507:32]
  reg [33:0] PMDU1_bits_Pctrl_mulres17_0; // @[SIMDU.scala 507:32]
  reg [33:0] PMDU1_bits_Pctrl_mulres17_1; // @[SIMDU.scala 507:32]
  reg [65:0] PMDU1_bits_Pctrl_mulres33_0; // @[SIMDU.scala 507:32]
  reg [129:0] PMDU1_bits_Pctrl_mulres65_0; // @[SIMDU.scala 507:32]
  reg  PMDU1_valid; // @[SIMDU.scala 509:28]
  wire  _GEN_3 = PMDU1_io_FirstStageFire ? 1'h0 : PMDU1_valid; // @[SIMDU.scala 511:19 512:{32,50}]
  wire  _T_12 = io_DecodeIn_0_InstNo <= io_DecodeIn_1_InstNo & io_DecodeIn_0_InstFlag == io_DecodeIn_1_InstFlag |
    io_DecodeIn_0_InstNo > io_DecodeIn_1_InstNo & io_DecodeIn_0_InstFlag != io_DecodeIn_1_InstFlag; // @[SIMDU.scala 450:101]
  wire  _T_13 = _T_12 ? 1'h0 : 1'h1; // @[SIMDU.scala 516:59]
  wire  firstidx = io_in_0_valid ? io_in_1_valid & _T_13 : 1'h1; // @[SIMDU.scala 516:21]
  wire  secondidx = ~firstidx; // @[SIMDU.scala 517:32]
  wire [4:0] _GEN_5 = firstidx ? io_DecodeIn_1_cf_instrType : io_DecodeIn_0_cf_instrType; // @[SIMDU.scala 518:{69,69}]
  wire  _GEN_7 = firstidx ? io_in_1_valid : io_in_0_valid; // @[SIMDU.scala 518:{30,30}]
  wire  _GEN_9 = firstidx ? io_DecodeIn_1_InstFlag : io_DecodeIn_0_InstFlag; // @[SIMDU.scala 522:{32,32}]
  wire [4:0] _GEN_11 = firstidx ? io_DecodeIn_1_InstNo : io_DecodeIn_0_InstNo; // @[SIMDU.scala 522:{32,32}]
  wire [63:0] _GEN_17 = firstidx ? io_DecodeIn_1_data_src3 : io_DecodeIn_0_data_src3; // @[SIMDU.scala 522:{32,32}]
  wire [63:0] _GEN_19 = firstidx ? io_DecodeIn_1_data_src2 : io_DecodeIn_0_data_src2; // @[SIMDU.scala 522:{32,32}]
  wire [63:0] _GEN_21 = firstidx ? io_DecodeIn_1_data_src1 : io_DecodeIn_0_data_src1; // @[SIMDU.scala 522:{32,32}]
  wire [4:0] _GEN_37 = firstidx ? io_DecodeIn_1_ctrl_rfDest : io_DecodeIn_0_ctrl_rfDest; // @[SIMDU.scala 522:{32,32}]
  wire  _GEN_39 = firstidx ? io_DecodeIn_1_ctrl_rfWen : io_DecodeIn_0_ctrl_rfWen; // @[SIMDU.scala 522:{32,32}]
  wire  _GEN_49 = firstidx ? io_DecodeIn_1_ctrl_func24 : io_DecodeIn_0_ctrl_func24; // @[SIMDU.scala 522:{32,32}]
  wire [2:0] _GEN_51 = firstidx ? io_DecodeIn_1_ctrl_funct3 : io_DecodeIn_0_ctrl_funct3; // @[SIMDU.scala 522:{32,32}]
  wire [6:0] _GEN_53 = firstidx ? io_DecodeIn_1_ctrl_fuOpType : io_DecodeIn_0_ctrl_fuOpType; // @[SIMDU.scala 522:{32,32}]
  wire [63:0] _GEN_63 = firstidx ? io_DecodeIn_1_cf_runahead_checkpoint_id : io_DecodeIn_0_cf_runahead_checkpoint_id; // @[SIMDU.scala 522:{32,32}]
  wire [38:0] _GEN_135 = firstidx ? io_DecodeIn_1_cf_pc : io_DecodeIn_0_cf_pc; // @[SIMDU.scala 522:{32,32}]
  wire  _T_23_isAdd_64 = secondidx ? PIDU0_io_Pctrl_isAdd_64 : PIDU1_io_Pctrl_isAdd_64; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdd_32 = secondidx ? PIDU0_io_Pctrl_isAdd_32 : PIDU1_io_Pctrl_isAdd_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdd_16 = secondidx ? PIDU0_io_Pctrl_isAdd_16 : PIDU1_io_Pctrl_isAdd_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdd_8 = secondidx ? PIDU0_io_Pctrl_isAdd_8 : PIDU1_io_Pctrl_isAdd_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdd_Q15 = secondidx ? PIDU0_io_Pctrl_isAdd_Q15 : PIDU1_io_Pctrl_isAdd_Q15; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdd_Q31 = secondidx ? PIDU0_io_Pctrl_isAdd_Q31 : PIDU1_io_Pctrl_isAdd_Q31; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdd_C31 = secondidx ? PIDU0_io_Pctrl_isAdd_C31 : PIDU1_io_Pctrl_isAdd_C31; // @[SIMDU.scala 523:38]
  wire  _T_23_isAve = secondidx ? PIDU0_io_Pctrl_isAve : PIDU1_io_Pctrl_isAve; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_64 = secondidx ? PIDU0_io_Pctrl_isSub_64 : PIDU1_io_Pctrl_isSub_64; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_32 = secondidx ? PIDU0_io_Pctrl_isSub_32 : PIDU1_io_Pctrl_isSub_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_16 = secondidx ? PIDU0_io_Pctrl_isSub_16 : PIDU1_io_Pctrl_isSub_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_8 = secondidx ? PIDU0_io_Pctrl_isSub_8 : PIDU1_io_Pctrl_isSub_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_Q15 = secondidx ? PIDU0_io_Pctrl_isSub_Q15 : PIDU1_io_Pctrl_isSub_Q15; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_Q31 = secondidx ? PIDU0_io_Pctrl_isSub_Q31 : PIDU1_io_Pctrl_isSub_Q31; // @[SIMDU.scala 523:38]
  wire  _T_23_isSub_C31 = secondidx ? PIDU0_io_Pctrl_isSub_C31 : PIDU1_io_Pctrl_isSub_C31; // @[SIMDU.scala 523:38]
  wire  _T_23_isCras_16 = secondidx ? PIDU0_io_Pctrl_isCras_16 : PIDU1_io_Pctrl_isCras_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isCrsa_16 = secondidx ? PIDU0_io_Pctrl_isCrsa_16 : PIDU1_io_Pctrl_isCrsa_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isCras_32 = secondidx ? PIDU0_io_Pctrl_isCras_32 : PIDU1_io_Pctrl_isCras_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isCrsa_32 = secondidx ? PIDU0_io_Pctrl_isCrsa_32 : PIDU1_io_Pctrl_isCrsa_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isStas_16 = secondidx ? PIDU0_io_Pctrl_isStas_16 : PIDU1_io_Pctrl_isStas_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isStsa_16 = secondidx ? PIDU0_io_Pctrl_isStsa_16 : PIDU1_io_Pctrl_isStsa_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isStas_32 = secondidx ? PIDU0_io_Pctrl_isStas_32 : PIDU1_io_Pctrl_isStas_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isStsa_32 = secondidx ? PIDU0_io_Pctrl_isStsa_32 : PIDU1_io_Pctrl_isStsa_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isComp_16 = secondidx ? PIDU0_io_Pctrl_isComp_16 : PIDU1_io_Pctrl_isComp_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isComp_8 = secondidx ? PIDU0_io_Pctrl_isComp_8 : PIDU1_io_Pctrl_isComp_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isCompare = secondidx ? PIDU0_io_Pctrl_isCompare : PIDU1_io_Pctrl_isCompare; // @[SIMDU.scala 523:38]
  wire  _T_23_isMaxMin_16 = secondidx ? PIDU0_io_Pctrl_isMaxMin_16 : PIDU1_io_Pctrl_isMaxMin_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isMaxMin_8 = secondidx ? PIDU0_io_Pctrl_isMaxMin_8 : PIDU1_io_Pctrl_isMaxMin_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isMaxMin_XLEN = secondidx ? PIDU0_io_Pctrl_isMaxMin_XLEN : PIDU1_io_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 523:38]
  wire  _T_23_isMaxMin_32 = secondidx ? PIDU0_io_Pctrl_isMaxMin_32 : PIDU1_io_Pctrl_isMaxMin_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isMaxMin = secondidx ? PIDU0_io_Pctrl_isMaxMin : PIDU1_io_Pctrl_isMaxMin; // @[SIMDU.scala 523:38]
  wire  _T_23_isPbs = secondidx ? PIDU0_io_Pctrl_isPbs : PIDU1_io_Pctrl_isPbs; // @[SIMDU.scala 523:38]
  wire  _T_23_isRs_16 = secondidx ? PIDU0_io_Pctrl_isRs_16 : PIDU1_io_Pctrl_isRs_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isLs_16 = secondidx ? PIDU0_io_Pctrl_isLs_16 : PIDU1_io_Pctrl_isLs_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isLR_16 = secondidx ? PIDU0_io_Pctrl_isLR_16 : PIDU1_io_Pctrl_isLR_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isRs_8 = secondidx ? PIDU0_io_Pctrl_isRs_8 : PIDU1_io_Pctrl_isRs_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isLs_8 = secondidx ? PIDU0_io_Pctrl_isLs_8 : PIDU1_io_Pctrl_isLs_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isLR_8 = secondidx ? PIDU0_io_Pctrl_isLR_8 : PIDU1_io_Pctrl_isLR_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isRs_32 = secondidx ? PIDU0_io_Pctrl_isRs_32 : PIDU1_io_Pctrl_isRs_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isLs_32 = secondidx ? PIDU0_io_Pctrl_isLs_32 : PIDU1_io_Pctrl_isLs_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isLR_32 = secondidx ? PIDU0_io_Pctrl_isLR_32 : PIDU1_io_Pctrl_isLR_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isLR_Q31 = secondidx ? PIDU0_io_Pctrl_isLR_Q31 : PIDU1_io_Pctrl_isLR_Q31; // @[SIMDU.scala 523:38]
  wire  _T_23_isLs_Q31 = secondidx ? PIDU0_io_Pctrl_isLs_Q31 : PIDU1_io_Pctrl_isLs_Q31; // @[SIMDU.scala 523:38]
  wire  _T_23_isRs_XLEN = secondidx ? PIDU0_io_Pctrl_isRs_XLEN : PIDU1_io_Pctrl_isRs_XLEN; // @[SIMDU.scala 523:38]
  wire  _T_23_isSRAIWU = secondidx ? PIDU0_io_Pctrl_isSRAIWU : PIDU1_io_Pctrl_isSRAIWU; // @[SIMDU.scala 523:38]
  wire  _T_23_isFSRW = secondidx ? PIDU0_io_Pctrl_isFSRW : PIDU1_io_Pctrl_isFSRW; // @[SIMDU.scala 523:38]
  wire  _T_23_isWext = secondidx ? PIDU0_io_Pctrl_isWext : PIDU1_io_Pctrl_isWext; // @[SIMDU.scala 523:38]
  wire  _T_23_isShifter = secondidx ? PIDU0_io_Pctrl_isShifter : PIDU1_io_Pctrl_isShifter; // @[SIMDU.scala 523:38]
  wire  _T_23_isClip_16 = secondidx ? PIDU0_io_Pctrl_isClip_16 : PIDU1_io_Pctrl_isClip_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isClip_8 = secondidx ? PIDU0_io_Pctrl_isClip_8 : PIDU1_io_Pctrl_isClip_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isclip_32 = secondidx ? PIDU0_io_Pctrl_isclip_32 : PIDU1_io_Pctrl_isclip_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isClip = secondidx ? PIDU0_io_Pctrl_isClip : PIDU1_io_Pctrl_isClip; // @[SIMDU.scala 523:38]
  wire  _T_23_isSat_16 = secondidx ? PIDU0_io_Pctrl_isSat_16 : PIDU1_io_Pctrl_isSat_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isSat_8 = secondidx ? PIDU0_io_Pctrl_isSat_8 : PIDU1_io_Pctrl_isSat_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isSat_32 = secondidx ? PIDU0_io_Pctrl_isSat_32 : PIDU1_io_Pctrl_isSat_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isSat_W = secondidx ? PIDU0_io_Pctrl_isSat_W : PIDU1_io_Pctrl_isSat_W; // @[SIMDU.scala 523:38]
  wire  _T_23_isSat = secondidx ? PIDU0_io_Pctrl_isSat : PIDU1_io_Pctrl_isSat; // @[SIMDU.scala 523:38]
  wire  _T_23_isCnt_16 = secondidx ? PIDU0_io_Pctrl_isCnt_16 : PIDU1_io_Pctrl_isCnt_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isCnt_8 = secondidx ? PIDU0_io_Pctrl_isCnt_8 : PIDU1_io_Pctrl_isCnt_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isCnt_32 = secondidx ? PIDU0_io_Pctrl_isCnt_32 : PIDU1_io_Pctrl_isCnt_32; // @[SIMDU.scala 523:38]
  wire  _T_23_isCnt = secondidx ? PIDU0_io_Pctrl_isCnt : PIDU1_io_Pctrl_isCnt; // @[SIMDU.scala 523:38]
  wire  _T_23_isSwap_16 = secondidx ? PIDU0_io_Pctrl_isSwap_16 : PIDU1_io_Pctrl_isSwap_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isSwap_8 = secondidx ? PIDU0_io_Pctrl_isSwap_8 : PIDU1_io_Pctrl_isSwap_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isSwap = secondidx ? PIDU0_io_Pctrl_isSwap : PIDU1_io_Pctrl_isSwap; // @[SIMDU.scala 523:38]
  wire  _T_23_isUnpack = secondidx ? PIDU0_io_Pctrl_isUnpack : PIDU1_io_Pctrl_isUnpack; // @[SIMDU.scala 523:38]
  wire  _T_23_isBitrev = secondidx ? PIDU0_io_Pctrl_isBitrev : PIDU1_io_Pctrl_isBitrev; // @[SIMDU.scala 523:38]
  wire  _T_23_isCmix = secondidx ? PIDU0_io_Pctrl_isCmix : PIDU1_io_Pctrl_isCmix; // @[SIMDU.scala 523:38]
  wire  _T_23_isInsertb = secondidx ? PIDU0_io_Pctrl_isInsertb : PIDU1_io_Pctrl_isInsertb; // @[SIMDU.scala 523:38]
  wire  _T_23_isPackbb = secondidx ? PIDU0_io_Pctrl_isPackbb : PIDU1_io_Pctrl_isPackbb; // @[SIMDU.scala 523:38]
  wire  _T_23_isPackbt = secondidx ? PIDU0_io_Pctrl_isPackbt : PIDU1_io_Pctrl_isPackbt; // @[SIMDU.scala 523:38]
  wire  _T_23_isPacktb = secondidx ? PIDU0_io_Pctrl_isPacktb : PIDU1_io_Pctrl_isPacktb; // @[SIMDU.scala 523:38]
  wire  _T_23_isPacktt = secondidx ? PIDU0_io_Pctrl_isPacktt : PIDU1_io_Pctrl_isPacktt; // @[SIMDU.scala 523:38]
  wire  _T_23_isPack = secondidx ? PIDU0_io_Pctrl_isPack : PIDU1_io_Pctrl_isPack; // @[SIMDU.scala 523:38]
  wire [7:0] _T_23_isSub = secondidx ? PIDU0_io_Pctrl_isSub : PIDU1_io_Pctrl_isSub; // @[SIMDU.scala 523:38]
  wire  _T_23_isAdder = secondidx ? PIDU0_io_Pctrl_isAdder : PIDU1_io_Pctrl_isAdder; // @[SIMDU.scala 523:38]
  wire  _T_23_SrcSigned = secondidx ? PIDU0_io_Pctrl_SrcSigned : PIDU1_io_Pctrl_SrcSigned; // @[SIMDU.scala 523:38]
  wire  _T_23_Saturating = secondidx ? PIDU0_io_Pctrl_Saturating : PIDU1_io_Pctrl_Saturating; // @[SIMDU.scala 523:38]
  wire  _T_23_Translation = secondidx ? PIDU0_io_Pctrl_Translation : PIDU1_io_Pctrl_Translation; // @[SIMDU.scala 523:38]
  wire  _T_23_LessEqual = secondidx ? PIDU0_io_Pctrl_LessEqual : PIDU1_io_Pctrl_LessEqual; // @[SIMDU.scala 523:38]
  wire  _T_23_LessThan = secondidx ? PIDU0_io_Pctrl_LessThan : PIDU1_io_Pctrl_LessThan; // @[SIMDU.scala 523:38]
  wire [79:0] _T_23_adderRes_ori = secondidx ? PIDU0_io_Pctrl_adderRes_ori : PIDU1_io_Pctrl_adderRes_ori; // @[SIMDU.scala 523:38]
  wire [63:0] _T_23_adderRes = secondidx ? PIDU0_io_Pctrl_adderRes : PIDU1_io_Pctrl_adderRes; // @[SIMDU.scala 523:38]
  wire [79:0] _T_23_adderRes_ori_drophighestbit = secondidx ? PIDU0_io_Pctrl_adderRes_ori_drophighestbit :
    PIDU1_io_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 523:38]
  wire  _T_23_Round = secondidx ? PIDU0_io_Pctrl_Round : PIDU1_io_Pctrl_Round; // @[SIMDU.scala 523:38]
  wire  _T_23_ShiftSigned = secondidx ? PIDU0_io_Pctrl_ShiftSigned : PIDU1_io_Pctrl_ShiftSigned; // @[SIMDU.scala 523:38]
  wire  _T_23_Arithmetic = secondidx ? PIDU0_io_Pctrl_Arithmetic : PIDU1_io_Pctrl_Arithmetic; // @[SIMDU.scala 523:38]
  wire  _T_23_isMul_16 = secondidx ? PIDU0_io_Pctrl_isMul_16 : PIDU1_io_Pctrl_isMul_16; // @[SIMDU.scala 523:38]
  wire  _T_23_isMul_8 = secondidx ? PIDU0_io_Pctrl_isMul_8 : PIDU1_io_Pctrl_isMul_8; // @[SIMDU.scala 523:38]
  wire  _T_23_isMSW_3232 = secondidx ? PIDU0_io_Pctrl_isMSW_3232 : PIDU1_io_Pctrl_isMSW_3232; // @[SIMDU.scala 523:38]
  wire  _T_23_isMSW_3216 = secondidx ? PIDU0_io_Pctrl_isMSW_3216 : PIDU1_io_Pctrl_isMSW_3216; // @[SIMDU.scala 523:38]
  wire  _T_23_isS1632 = secondidx ? PIDU0_io_Pctrl_isS1632 : PIDU1_io_Pctrl_isS1632; // @[SIMDU.scala 523:38]
  wire  _T_23_isS1664 = secondidx ? PIDU0_io_Pctrl_isS1664 : PIDU1_io_Pctrl_isS1664; // @[SIMDU.scala 523:38]
  wire  _T_23_is832 = secondidx ? PIDU0_io_Pctrl_is832 : PIDU1_io_Pctrl_is832; // @[SIMDU.scala 523:38]
  wire  _T_23_is3264 = secondidx ? PIDU0_io_Pctrl_is3264 : PIDU1_io_Pctrl_is3264; // @[SIMDU.scala 523:38]
  wire  _T_23_is1664 = secondidx ? PIDU0_io_Pctrl_is1664 : PIDU1_io_Pctrl_is1664; // @[SIMDU.scala 523:38]
  wire  _T_23_isQ15orQ31 = secondidx ? PIDU0_io_Pctrl_isQ15orQ31 : PIDU1_io_Pctrl_isQ15orQ31; // @[SIMDU.scala 523:38]
  wire  _T_23_isC31 = secondidx ? PIDU0_io_Pctrl_isC31 : PIDU1_io_Pctrl_isC31; // @[SIMDU.scala 523:38]
  wire  _T_23_isQ15_64ONLY = secondidx ? PIDU0_io_Pctrl_isQ15_64ONLY : PIDU1_io_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 523:38]
  wire  _T_23_isQ63_64ONLY = secondidx ? PIDU0_io_Pctrl_isQ63_64ONLY : PIDU1_io_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 523:38]
  wire  _T_23_isMul_32_64ONLY = secondidx ? PIDU0_io_Pctrl_isMul_32_64ONLY : PIDU1_io_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 523:38]
  wire  _T_23_isPMA_64ONLY = secondidx ? PIDU0_io_Pctrl_isPMA_64ONLY : PIDU1_io_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 523:38]
  wire [17:0] _T_23_mulres9_0 = secondidx ? PIDU0_io_Pctrl_mulres9_0 : PIDU1_io_Pctrl_mulres9_0; // @[SIMDU.scala 523:38]
  wire [17:0] _T_23_mulres9_1 = secondidx ? PIDU0_io_Pctrl_mulres9_1 : PIDU1_io_Pctrl_mulres9_1; // @[SIMDU.scala 523:38]
  wire [17:0] _T_23_mulres9_2 = secondidx ? PIDU0_io_Pctrl_mulres9_2 : PIDU1_io_Pctrl_mulres9_2; // @[SIMDU.scala 523:38]
  wire [17:0] _T_23_mulres9_3 = secondidx ? PIDU0_io_Pctrl_mulres9_3 : PIDU1_io_Pctrl_mulres9_3; // @[SIMDU.scala 523:38]
  wire [33:0] _T_23_mulres17_0 = secondidx ? PIDU0_io_Pctrl_mulres17_0 : PIDU1_io_Pctrl_mulres17_0; // @[SIMDU.scala 523:38]
  wire [33:0] _T_23_mulres17_1 = secondidx ? PIDU0_io_Pctrl_mulres17_1 : PIDU1_io_Pctrl_mulres17_1; // @[SIMDU.scala 523:38]
  wire [65:0] _T_23_mulres33_0 = secondidx ? PIDU0_io_Pctrl_mulres33_0 : PIDU1_io_Pctrl_mulres33_0; // @[SIMDU.scala 523:38]
  wire [129:0] _T_23_mulres65_0 = secondidx ? PIDU0_io_Pctrl_mulres65_0 : PIDU1_io_Pctrl_mulres65_0; // @[SIMDU.scala 523:38]
  wire  _GEN_142 = PALU1_io_in_ready; // @[SIMDU.scala 525:34 526:25]
  wire  _GEN_143 = PALU1_io_in_ready | _GEN_1; // @[SIMDU.scala 525:34 527:24]
  wire  _GEN_144 = PALU1_io_in_ready ? _GEN_9 : PALU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [4:0] _GEN_145 = PALU1_io_in_ready ? _GEN_11 : PALU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [63:0] _GEN_148 = PALU1_io_in_ready ? _GEN_17 : PALU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [63:0] _GEN_149 = PALU1_io_in_ready ? _GEN_19 : PALU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [63:0] _GEN_150 = PALU1_io_in_ready ? _GEN_21 : PALU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [4:0] _GEN_158 = PALU1_io_in_ready ? _GEN_37 : PALU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 491:19 525:34 528:32]
  wire  _GEN_159 = PALU1_io_in_ready ? _GEN_39 : PALU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 491:19 525:34 528:32]
  wire  _GEN_164 = PALU1_io_in_ready ? _GEN_49 : PALU1_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [2:0] _GEN_165 = PALU1_io_in_ready ? _GEN_51 : PALU1_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [6:0] _GEN_166 = PALU1_io_in_ready ? _GEN_53 : PALU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [63:0] _GEN_172 = PALU1_io_in_ready ? _GEN_63 : PALU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 491:19 525:34 528:32]
  wire [38:0] _GEN_208 = PALU1_io_in_ready ? _GEN_135 : PALU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 491:19 525:34 528:32]
  wire  _GEN_233 = PALU1_io_in_ready ? _T_23_Arithmetic : PALU1_bits_Pctrl_Arithmetic; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_234 = PALU1_io_in_ready ? _T_23_ShiftSigned : PALU1_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_235 = PALU1_io_in_ready ? _T_23_Round : PALU1_bits_Pctrl_Round; // @[SIMDU.scala 491:19 525:34 529:32]
  wire [79:0] _GEN_236 = PALU1_io_in_ready ? _T_23_adderRes_ori_drophighestbit :
    PALU1_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 491:19 525:34 529:32]
  wire [63:0] _GEN_237 = PALU1_io_in_ready ? _T_23_adderRes : PALU1_bits_Pctrl_adderRes; // @[SIMDU.scala 491:19 525:34 529:32]
  wire [79:0] _GEN_238 = PALU1_io_in_ready ? _T_23_adderRes_ori : PALU1_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_239 = PALU1_io_in_ready ? _T_23_LessThan : PALU1_bits_Pctrl_LessThan; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_240 = PALU1_io_in_ready ? _T_23_LessEqual : PALU1_bits_Pctrl_LessEqual; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_241 = PALU1_io_in_ready ? _T_23_Translation : PALU1_bits_Pctrl_Translation; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_242 = PALU1_io_in_ready ? _T_23_Saturating : PALU1_bits_Pctrl_Saturating; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_243 = PALU1_io_in_ready ? _T_23_SrcSigned : PALU1_bits_Pctrl_SrcSigned; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_244 = PALU1_io_in_ready ? _T_23_isAdder : PALU1_bits_Pctrl_isAdder; // @[SIMDU.scala 491:19 525:34 529:32]
  wire [7:0] _GEN_245 = PALU1_io_in_ready ? _T_23_isSub : PALU1_bits_Pctrl_isSub; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_246 = PALU1_io_in_ready ? _T_23_isPack : PALU1_bits_Pctrl_isPack; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_247 = PALU1_io_in_ready ? _T_23_isPacktt : PALU1_bits_Pctrl_isPacktt; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_248 = PALU1_io_in_ready ? _T_23_isPacktb : PALU1_bits_Pctrl_isPacktb; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_249 = PALU1_io_in_ready ? _T_23_isPackbt : PALU1_bits_Pctrl_isPackbt; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_250 = PALU1_io_in_ready ? _T_23_isPackbb : PALU1_bits_Pctrl_isPackbb; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_251 = PALU1_io_in_ready ? _T_23_isInsertb : PALU1_bits_Pctrl_isInsertb; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_252 = PALU1_io_in_ready ? _T_23_isCmix : PALU1_bits_Pctrl_isCmix; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_253 = PALU1_io_in_ready ? _T_23_isBitrev : PALU1_bits_Pctrl_isBitrev; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_254 = PALU1_io_in_ready ? _T_23_isUnpack : PALU1_bits_Pctrl_isUnpack; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_255 = PALU1_io_in_ready ? _T_23_isSwap : PALU1_bits_Pctrl_isSwap; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_256 = PALU1_io_in_ready ? _T_23_isSwap_8 : PALU1_bits_Pctrl_isSwap_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_257 = PALU1_io_in_ready ? _T_23_isSwap_16 : PALU1_bits_Pctrl_isSwap_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_258 = PALU1_io_in_ready ? _T_23_isCnt : PALU1_bits_Pctrl_isCnt; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_259 = PALU1_io_in_ready ? _T_23_isCnt_32 : PALU1_bits_Pctrl_isCnt_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_260 = PALU1_io_in_ready ? _T_23_isCnt_8 : PALU1_bits_Pctrl_isCnt_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_261 = PALU1_io_in_ready ? _T_23_isCnt_16 : PALU1_bits_Pctrl_isCnt_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_262 = PALU1_io_in_ready ? _T_23_isSat : PALU1_bits_Pctrl_isSat; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_263 = PALU1_io_in_ready ? _T_23_isSat_W : PALU1_bits_Pctrl_isSat_W; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_264 = PALU1_io_in_ready ? _T_23_isSat_32 : PALU1_bits_Pctrl_isSat_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_265 = PALU1_io_in_ready ? _T_23_isSat_8 : PALU1_bits_Pctrl_isSat_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_266 = PALU1_io_in_ready ? _T_23_isSat_16 : PALU1_bits_Pctrl_isSat_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_267 = PALU1_io_in_ready ? _T_23_isClip : PALU1_bits_Pctrl_isClip; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_268 = PALU1_io_in_ready ? _T_23_isclip_32 : PALU1_bits_Pctrl_isclip_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_269 = PALU1_io_in_ready ? _T_23_isClip_8 : PALU1_bits_Pctrl_isClip_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_270 = PALU1_io_in_ready ? _T_23_isClip_16 : PALU1_bits_Pctrl_isClip_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_271 = PALU1_io_in_ready ? _T_23_isShifter : PALU1_bits_Pctrl_isShifter; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_272 = PALU1_io_in_ready ? _T_23_isWext : PALU1_bits_Pctrl_isWext; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_273 = PALU1_io_in_ready ? _T_23_isFSRW : PALU1_bits_Pctrl_isFSRW; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_274 = PALU1_io_in_ready ? _T_23_isSRAIWU : PALU1_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_275 = PALU1_io_in_ready ? _T_23_isRs_XLEN : PALU1_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_276 = PALU1_io_in_ready ? _T_23_isLs_Q31 : PALU1_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_277 = PALU1_io_in_ready ? _T_23_isLR_Q31 : PALU1_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_278 = PALU1_io_in_ready ? _T_23_isLR_32 : PALU1_bits_Pctrl_isLR_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_279 = PALU1_io_in_ready ? _T_23_isLs_32 : PALU1_bits_Pctrl_isLs_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_280 = PALU1_io_in_ready ? _T_23_isRs_32 : PALU1_bits_Pctrl_isRs_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_281 = PALU1_io_in_ready ? _T_23_isLR_8 : PALU1_bits_Pctrl_isLR_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_282 = PALU1_io_in_ready ? _T_23_isLs_8 : PALU1_bits_Pctrl_isLs_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_283 = PALU1_io_in_ready ? _T_23_isRs_8 : PALU1_bits_Pctrl_isRs_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_284 = PALU1_io_in_ready ? _T_23_isLR_16 : PALU1_bits_Pctrl_isLR_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_285 = PALU1_io_in_ready ? _T_23_isLs_16 : PALU1_bits_Pctrl_isLs_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_286 = PALU1_io_in_ready ? _T_23_isRs_16 : PALU1_bits_Pctrl_isRs_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_287 = PALU1_io_in_ready ? _T_23_isPbs : PALU1_bits_Pctrl_isPbs; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_288 = PALU1_io_in_ready ? _T_23_isMaxMin : PALU1_bits_Pctrl_isMaxMin; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_289 = PALU1_io_in_ready ? _T_23_isMaxMin_32 : PALU1_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_290 = PALU1_io_in_ready ? _T_23_isMaxMin_XLEN : PALU1_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_291 = PALU1_io_in_ready ? _T_23_isMaxMin_8 : PALU1_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_292 = PALU1_io_in_ready ? _T_23_isMaxMin_16 : PALU1_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_293 = PALU1_io_in_ready ? _T_23_isCompare : PALU1_bits_Pctrl_isCompare; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_294 = PALU1_io_in_ready ? _T_23_isComp_8 : PALU1_bits_Pctrl_isComp_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_295 = PALU1_io_in_ready ? _T_23_isComp_16 : PALU1_bits_Pctrl_isComp_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_297 = PALU1_io_in_ready ? _T_23_isStsa_32 : PALU1_bits_Pctrl_isStsa_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_298 = PALU1_io_in_ready ? _T_23_isStas_32 : PALU1_bits_Pctrl_isStas_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_299 = PALU1_io_in_ready ? _T_23_isStsa_16 : PALU1_bits_Pctrl_isStsa_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_300 = PALU1_io_in_ready ? _T_23_isStas_16 : PALU1_bits_Pctrl_isStas_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_302 = PALU1_io_in_ready ? _T_23_isCrsa_32 : PALU1_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_303 = PALU1_io_in_ready ? _T_23_isCras_32 : PALU1_bits_Pctrl_isCras_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_304 = PALU1_io_in_ready ? _T_23_isCrsa_16 : PALU1_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_305 = PALU1_io_in_ready ? _T_23_isCras_16 : PALU1_bits_Pctrl_isCras_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_306 = PALU1_io_in_ready ? _T_23_isSub_C31 : PALU1_bits_Pctrl_isSub_C31; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_307 = PALU1_io_in_ready ? _T_23_isSub_Q31 : PALU1_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_308 = PALU1_io_in_ready ? _T_23_isSub_Q15 : PALU1_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_309 = PALU1_io_in_ready ? _T_23_isSub_8 : PALU1_bits_Pctrl_isSub_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_310 = PALU1_io_in_ready ? _T_23_isSub_16 : PALU1_bits_Pctrl_isSub_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_311 = PALU1_io_in_ready ? _T_23_isSub_32 : PALU1_bits_Pctrl_isSub_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_312 = PALU1_io_in_ready ? _T_23_isSub_64 : PALU1_bits_Pctrl_isSub_64; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_314 = PALU1_io_in_ready ? _T_23_isAve : PALU1_bits_Pctrl_isAve; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_315 = PALU1_io_in_ready ? _T_23_isAdd_C31 : PALU1_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_316 = PALU1_io_in_ready ? _T_23_isAdd_Q31 : PALU1_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_317 = PALU1_io_in_ready ? _T_23_isAdd_Q15 : PALU1_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_318 = PALU1_io_in_ready ? _T_23_isAdd_8 : PALU1_bits_Pctrl_isAdd_8; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_319 = PALU1_io_in_ready ? _T_23_isAdd_16 : PALU1_bits_Pctrl_isAdd_16; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_320 = PALU1_io_in_ready ? _T_23_isAdd_32 : PALU1_bits_Pctrl_isAdd_32; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_321 = PALU1_io_in_ready ? _T_23_isAdd_64 : PALU1_bits_Pctrl_isAdd_64; // @[SIMDU.scala 491:19 525:34 529:32]
  wire  _GEN_322 = PALU1_io_in_ready & secondidx; // @[SIMDU.scala 472:24 525:34]
  wire  _GEN_323 = PALU1_io_in_ready & firstidx; // @[SIMDU.scala 473:24 525:34]
  wire  _GEN_324 = PALU0_io_in_ready; // @[SIMDU.scala 519:28 520:25]
  wire  _GEN_325 = PALU0_io_in_ready | _GEN_0; // @[SIMDU.scala 519:28 521:24]
  wire  _GEN_326 = PALU0_io_in_ready ? _GEN_9 : PALU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [4:0] _GEN_327 = PALU0_io_in_ready ? _GEN_11 : PALU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [63:0] _GEN_330 = PALU0_io_in_ready ? _GEN_17 : PALU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [63:0] _GEN_331 = PALU0_io_in_ready ? _GEN_19 : PALU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [63:0] _GEN_332 = PALU0_io_in_ready ? _GEN_21 : PALU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [4:0] _GEN_340 = PALU0_io_in_ready ? _GEN_37 : PALU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 483:19 519:28 522:32]
  wire  _GEN_341 = PALU0_io_in_ready ? _GEN_39 : PALU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 483:19 519:28 522:32]
  wire  _GEN_346 = PALU0_io_in_ready ? _GEN_49 : PALU0_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [2:0] _GEN_347 = PALU0_io_in_ready ? _GEN_51 : PALU0_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [6:0] _GEN_348 = PALU0_io_in_ready ? _GEN_53 : PALU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [63:0] _GEN_354 = PALU0_io_in_ready ? _GEN_63 : PALU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 483:19 519:28 522:32]
  wire [38:0] _GEN_390 = PALU0_io_in_ready ? _GEN_135 : PALU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 483:19 519:28 522:32]
  wire  _GEN_415 = PALU0_io_in_ready ? _T_23_Arithmetic : PALU0_bits_Pctrl_Arithmetic; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_416 = PALU0_io_in_ready ? _T_23_ShiftSigned : PALU0_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_417 = PALU0_io_in_ready ? _T_23_Round : PALU0_bits_Pctrl_Round; // @[SIMDU.scala 483:19 519:28 523:32]
  wire [79:0] _GEN_418 = PALU0_io_in_ready ? _T_23_adderRes_ori_drophighestbit :
    PALU0_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 483:19 519:28 523:32]
  wire [63:0] _GEN_419 = PALU0_io_in_ready ? _T_23_adderRes : PALU0_bits_Pctrl_adderRes; // @[SIMDU.scala 483:19 519:28 523:32]
  wire [79:0] _GEN_420 = PALU0_io_in_ready ? _T_23_adderRes_ori : PALU0_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_421 = PALU0_io_in_ready ? _T_23_LessThan : PALU0_bits_Pctrl_LessThan; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_422 = PALU0_io_in_ready ? _T_23_LessEqual : PALU0_bits_Pctrl_LessEqual; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_423 = PALU0_io_in_ready ? _T_23_Translation : PALU0_bits_Pctrl_Translation; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_424 = PALU0_io_in_ready ? _T_23_Saturating : PALU0_bits_Pctrl_Saturating; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_425 = PALU0_io_in_ready ? _T_23_SrcSigned : PALU0_bits_Pctrl_SrcSigned; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_426 = PALU0_io_in_ready ? _T_23_isAdder : PALU0_bits_Pctrl_isAdder; // @[SIMDU.scala 483:19 519:28 523:32]
  wire [7:0] _GEN_427 = PALU0_io_in_ready ? _T_23_isSub : PALU0_bits_Pctrl_isSub; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_428 = PALU0_io_in_ready ? _T_23_isPack : PALU0_bits_Pctrl_isPack; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_429 = PALU0_io_in_ready ? _T_23_isPacktt : PALU0_bits_Pctrl_isPacktt; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_430 = PALU0_io_in_ready ? _T_23_isPacktb : PALU0_bits_Pctrl_isPacktb; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_431 = PALU0_io_in_ready ? _T_23_isPackbt : PALU0_bits_Pctrl_isPackbt; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_432 = PALU0_io_in_ready ? _T_23_isPackbb : PALU0_bits_Pctrl_isPackbb; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_433 = PALU0_io_in_ready ? _T_23_isInsertb : PALU0_bits_Pctrl_isInsertb; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_434 = PALU0_io_in_ready ? _T_23_isCmix : PALU0_bits_Pctrl_isCmix; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_435 = PALU0_io_in_ready ? _T_23_isBitrev : PALU0_bits_Pctrl_isBitrev; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_436 = PALU0_io_in_ready ? _T_23_isUnpack : PALU0_bits_Pctrl_isUnpack; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_437 = PALU0_io_in_ready ? _T_23_isSwap : PALU0_bits_Pctrl_isSwap; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_438 = PALU0_io_in_ready ? _T_23_isSwap_8 : PALU0_bits_Pctrl_isSwap_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_439 = PALU0_io_in_ready ? _T_23_isSwap_16 : PALU0_bits_Pctrl_isSwap_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_440 = PALU0_io_in_ready ? _T_23_isCnt : PALU0_bits_Pctrl_isCnt; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_441 = PALU0_io_in_ready ? _T_23_isCnt_32 : PALU0_bits_Pctrl_isCnt_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_442 = PALU0_io_in_ready ? _T_23_isCnt_8 : PALU0_bits_Pctrl_isCnt_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_443 = PALU0_io_in_ready ? _T_23_isCnt_16 : PALU0_bits_Pctrl_isCnt_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_444 = PALU0_io_in_ready ? _T_23_isSat : PALU0_bits_Pctrl_isSat; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_445 = PALU0_io_in_ready ? _T_23_isSat_W : PALU0_bits_Pctrl_isSat_W; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_446 = PALU0_io_in_ready ? _T_23_isSat_32 : PALU0_bits_Pctrl_isSat_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_447 = PALU0_io_in_ready ? _T_23_isSat_8 : PALU0_bits_Pctrl_isSat_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_448 = PALU0_io_in_ready ? _T_23_isSat_16 : PALU0_bits_Pctrl_isSat_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_449 = PALU0_io_in_ready ? _T_23_isClip : PALU0_bits_Pctrl_isClip; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_450 = PALU0_io_in_ready ? _T_23_isclip_32 : PALU0_bits_Pctrl_isclip_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_451 = PALU0_io_in_ready ? _T_23_isClip_8 : PALU0_bits_Pctrl_isClip_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_452 = PALU0_io_in_ready ? _T_23_isClip_16 : PALU0_bits_Pctrl_isClip_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_453 = PALU0_io_in_ready ? _T_23_isShifter : PALU0_bits_Pctrl_isShifter; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_454 = PALU0_io_in_ready ? _T_23_isWext : PALU0_bits_Pctrl_isWext; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_455 = PALU0_io_in_ready ? _T_23_isFSRW : PALU0_bits_Pctrl_isFSRW; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_456 = PALU0_io_in_ready ? _T_23_isSRAIWU : PALU0_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_457 = PALU0_io_in_ready ? _T_23_isRs_XLEN : PALU0_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_458 = PALU0_io_in_ready ? _T_23_isLs_Q31 : PALU0_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_459 = PALU0_io_in_ready ? _T_23_isLR_Q31 : PALU0_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_460 = PALU0_io_in_ready ? _T_23_isLR_32 : PALU0_bits_Pctrl_isLR_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_461 = PALU0_io_in_ready ? _T_23_isLs_32 : PALU0_bits_Pctrl_isLs_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_462 = PALU0_io_in_ready ? _T_23_isRs_32 : PALU0_bits_Pctrl_isRs_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_463 = PALU0_io_in_ready ? _T_23_isLR_8 : PALU0_bits_Pctrl_isLR_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_464 = PALU0_io_in_ready ? _T_23_isLs_8 : PALU0_bits_Pctrl_isLs_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_465 = PALU0_io_in_ready ? _T_23_isRs_8 : PALU0_bits_Pctrl_isRs_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_466 = PALU0_io_in_ready ? _T_23_isLR_16 : PALU0_bits_Pctrl_isLR_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_467 = PALU0_io_in_ready ? _T_23_isLs_16 : PALU0_bits_Pctrl_isLs_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_468 = PALU0_io_in_ready ? _T_23_isRs_16 : PALU0_bits_Pctrl_isRs_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_469 = PALU0_io_in_ready ? _T_23_isPbs : PALU0_bits_Pctrl_isPbs; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_470 = PALU0_io_in_ready ? _T_23_isMaxMin : PALU0_bits_Pctrl_isMaxMin; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_471 = PALU0_io_in_ready ? _T_23_isMaxMin_32 : PALU0_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_472 = PALU0_io_in_ready ? _T_23_isMaxMin_XLEN : PALU0_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_473 = PALU0_io_in_ready ? _T_23_isMaxMin_8 : PALU0_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_474 = PALU0_io_in_ready ? _T_23_isMaxMin_16 : PALU0_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_475 = PALU0_io_in_ready ? _T_23_isCompare : PALU0_bits_Pctrl_isCompare; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_476 = PALU0_io_in_ready ? _T_23_isComp_8 : PALU0_bits_Pctrl_isComp_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_477 = PALU0_io_in_ready ? _T_23_isComp_16 : PALU0_bits_Pctrl_isComp_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_479 = PALU0_io_in_ready ? _T_23_isStsa_32 : PALU0_bits_Pctrl_isStsa_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_480 = PALU0_io_in_ready ? _T_23_isStas_32 : PALU0_bits_Pctrl_isStas_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_481 = PALU0_io_in_ready ? _T_23_isStsa_16 : PALU0_bits_Pctrl_isStsa_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_482 = PALU0_io_in_ready ? _T_23_isStas_16 : PALU0_bits_Pctrl_isStas_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_484 = PALU0_io_in_ready ? _T_23_isCrsa_32 : PALU0_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_485 = PALU0_io_in_ready ? _T_23_isCras_32 : PALU0_bits_Pctrl_isCras_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_486 = PALU0_io_in_ready ? _T_23_isCrsa_16 : PALU0_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_487 = PALU0_io_in_ready ? _T_23_isCras_16 : PALU0_bits_Pctrl_isCras_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_488 = PALU0_io_in_ready ? _T_23_isSub_C31 : PALU0_bits_Pctrl_isSub_C31; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_489 = PALU0_io_in_ready ? _T_23_isSub_Q31 : PALU0_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_490 = PALU0_io_in_ready ? _T_23_isSub_Q15 : PALU0_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_491 = PALU0_io_in_ready ? _T_23_isSub_8 : PALU0_bits_Pctrl_isSub_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_492 = PALU0_io_in_ready ? _T_23_isSub_16 : PALU0_bits_Pctrl_isSub_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_493 = PALU0_io_in_ready ? _T_23_isSub_32 : PALU0_bits_Pctrl_isSub_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_494 = PALU0_io_in_ready ? _T_23_isSub_64 : PALU0_bits_Pctrl_isSub_64; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_496 = PALU0_io_in_ready ? _T_23_isAve : PALU0_bits_Pctrl_isAve; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_497 = PALU0_io_in_ready ? _T_23_isAdd_C31 : PALU0_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_498 = PALU0_io_in_ready ? _T_23_isAdd_Q31 : PALU0_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_499 = PALU0_io_in_ready ? _T_23_isAdd_Q15 : PALU0_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_500 = PALU0_io_in_ready ? _T_23_isAdd_8 : PALU0_bits_Pctrl_isAdd_8; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_501 = PALU0_io_in_ready ? _T_23_isAdd_16 : PALU0_bits_Pctrl_isAdd_16; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_502 = PALU0_io_in_ready ? _T_23_isAdd_32 : PALU0_bits_Pctrl_isAdd_32; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_503 = PALU0_io_in_ready ? _T_23_isAdd_64 : PALU0_bits_Pctrl_isAdd_64; // @[SIMDU.scala 483:19 519:28 523:32]
  wire  _GEN_504 = PALU0_io_in_ready ? secondidx : _GEN_322; // @[SIMDU.scala 519:28]
  wire  _GEN_505 = PALU0_io_in_ready ? firstidx : _GEN_323; // @[SIMDU.scala 519:28]
  wire  _GEN_506 = PALU0_io_in_ready ? 1'h0 : _GEN_142; // @[SIMDU.scala 519:28]
  wire  _GEN_507 = PALU0_io_in_ready ? _GEN_1 : _GEN_143; // @[SIMDU.scala 519:28]
  wire  _GEN_508 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_InstFlag : _GEN_144; // @[SIMDU.scala 491:19 519:28]
  wire [4:0] _GEN_509 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_InstNo : _GEN_145; // @[SIMDU.scala 491:19 519:28]
  wire [63:0] _GEN_512 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_data_src3 : _GEN_148; // @[SIMDU.scala 491:19 519:28]
  wire [63:0] _GEN_513 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_data_src2 : _GEN_149; // @[SIMDU.scala 491:19 519:28]
  wire [63:0] _GEN_514 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_data_src1 : _GEN_150; // @[SIMDU.scala 491:19 519:28]
  wire [4:0] _GEN_522 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_ctrl_rfDest : _GEN_158; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_523 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_ctrl_rfWen : _GEN_159; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_528 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_ctrl_func24 : _GEN_164; // @[SIMDU.scala 491:19 519:28]
  wire [2:0] _GEN_529 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_ctrl_funct3 : _GEN_165; // @[SIMDU.scala 491:19 519:28]
  wire [6:0] _GEN_530 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_ctrl_fuOpType : _GEN_166; // @[SIMDU.scala 491:19 519:28]
  wire [63:0] _GEN_536 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_cf_runahead_checkpoint_id : _GEN_172; // @[SIMDU.scala 491:19 519:28]
  wire [38:0] _GEN_572 = PALU0_io_in_ready ? PALU1_bits_DecodeIn_cf_pc : _GEN_208; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_597 = PALU0_io_in_ready ? PALU1_bits_Pctrl_Arithmetic : _GEN_233; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_598 = PALU0_io_in_ready ? PALU1_bits_Pctrl_ShiftSigned : _GEN_234; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_599 = PALU0_io_in_ready ? PALU1_bits_Pctrl_Round : _GEN_235; // @[SIMDU.scala 491:19 519:28]
  wire [79:0] _GEN_600 = PALU0_io_in_ready ? PALU1_bits_Pctrl_adderRes_ori_drophighestbit : _GEN_236; // @[SIMDU.scala 491:19 519:28]
  wire [63:0] _GEN_601 = PALU0_io_in_ready ? PALU1_bits_Pctrl_adderRes : _GEN_237; // @[SIMDU.scala 491:19 519:28]
  wire [79:0] _GEN_602 = PALU0_io_in_ready ? PALU1_bits_Pctrl_adderRes_ori : _GEN_238; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_603 = PALU0_io_in_ready ? PALU1_bits_Pctrl_LessThan : _GEN_239; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_604 = PALU0_io_in_ready ? PALU1_bits_Pctrl_LessEqual : _GEN_240; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_605 = PALU0_io_in_ready ? PALU1_bits_Pctrl_Translation : _GEN_241; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_606 = PALU0_io_in_ready ? PALU1_bits_Pctrl_Saturating : _GEN_242; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_607 = PALU0_io_in_ready ? PALU1_bits_Pctrl_SrcSigned : _GEN_243; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_608 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdder : _GEN_244; // @[SIMDU.scala 491:19 519:28]
  wire [7:0] _GEN_609 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub : _GEN_245; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_610 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isPack : _GEN_246; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_611 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isPacktt : _GEN_247; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_612 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isPacktb : _GEN_248; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_613 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isPackbt : _GEN_249; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_614 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isPackbb : _GEN_250; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_615 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isInsertb : _GEN_251; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_616 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCmix : _GEN_252; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_617 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isBitrev : _GEN_253; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_618 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isUnpack : _GEN_254; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_619 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSwap : _GEN_255; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_620 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSwap_8 : _GEN_256; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_621 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSwap_16 : _GEN_257; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_622 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCnt : _GEN_258; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_623 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCnt_32 : _GEN_259; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_624 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCnt_8 : _GEN_260; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_625 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCnt_16 : _GEN_261; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_626 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSat : _GEN_262; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_627 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSat_W : _GEN_263; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_628 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSat_32 : _GEN_264; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_629 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSat_8 : _GEN_265; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_630 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSat_16 : _GEN_266; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_631 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isClip : _GEN_267; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_632 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isclip_32 : _GEN_268; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_633 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isClip_8 : _GEN_269; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_634 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isClip_16 : _GEN_270; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_635 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isShifter : _GEN_271; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_636 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isWext : _GEN_272; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_637 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isFSRW : _GEN_273; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_638 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSRAIWU : _GEN_274; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_639 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isRs_XLEN : _GEN_275; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_640 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLs_Q31 : _GEN_276; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_641 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLR_Q31 : _GEN_277; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_642 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLR_32 : _GEN_278; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_643 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLs_32 : _GEN_279; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_644 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isRs_32 : _GEN_280; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_645 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLR_8 : _GEN_281; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_646 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLs_8 : _GEN_282; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_647 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isRs_8 : _GEN_283; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_648 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLR_16 : _GEN_284; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_649 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isLs_16 : _GEN_285; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_650 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isRs_16 : _GEN_286; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_651 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isPbs : _GEN_287; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_652 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isMaxMin : _GEN_288; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_653 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isMaxMin_32 : _GEN_289; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_654 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isMaxMin_XLEN : _GEN_290; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_655 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isMaxMin_8 : _GEN_291; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_656 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isMaxMin_16 : _GEN_292; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_657 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCompare : _GEN_293; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_658 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isComp_8 : _GEN_294; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_659 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isComp_16 : _GEN_295; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_661 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isStsa_32 : _GEN_297; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_662 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isStas_32 : _GEN_298; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_663 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isStsa_16 : _GEN_299; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_664 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isStas_16 : _GEN_300; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_666 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCrsa_32 : _GEN_302; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_667 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCras_32 : _GEN_303; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_668 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCrsa_16 : _GEN_304; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_669 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isCras_16 : _GEN_305; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_670 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_C31 : _GEN_306; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_671 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_Q31 : _GEN_307; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_672 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_Q15 : _GEN_308; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_673 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_8 : _GEN_309; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_674 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_16 : _GEN_310; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_675 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_32 : _GEN_311; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_676 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isSub_64 : _GEN_312; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_678 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAve : _GEN_314; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_679 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_C31 : _GEN_315; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_680 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_Q31 : _GEN_316; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_681 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_Q15 : _GEN_317; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_682 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_8 : _GEN_318; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_683 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_16 : _GEN_319; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_684 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_32 : _GEN_320; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_685 = PALU0_io_in_ready ? PALU1_bits_Pctrl_isAdd_64 : _GEN_321; // @[SIMDU.scala 491:19 519:28]
  wire  _GEN_690 = PMDU1_io_in_ready; // @[SIMDU.scala 539:34 540:25]
  wire  _GEN_691 = PMDU1_io_in_ready | _GEN_3; // @[SIMDU.scala 539:34 541:24]
  wire  _GEN_692 = PMDU1_io_in_ready ? _GEN_9 : PMDU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [4:0] _GEN_693 = PMDU1_io_in_ready ? _GEN_11 : PMDU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [63:0] _GEN_696 = PMDU1_io_in_ready ? _GEN_17 : PMDU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [63:0] _GEN_697 = PMDU1_io_in_ready ? _GEN_19 : PMDU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [63:0] _GEN_698 = PMDU1_io_in_ready ? _GEN_21 : PMDU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [4:0] _GEN_706 = PMDU1_io_in_ready ? _GEN_37 : PMDU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 508:19 539:34 542:32]
  wire  _GEN_707 = PMDU1_io_in_ready ? _GEN_39 : PMDU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [6:0] _GEN_714 = PMDU1_io_in_ready ? _GEN_53 : PMDU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [63:0] _GEN_720 = PMDU1_io_in_ready ? _GEN_63 : PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [38:0] _GEN_756 = PMDU1_io_in_ready ? _GEN_135 : PMDU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 508:19 539:34 542:32]
  wire [129:0] _GEN_758 = PMDU1_io_in_ready ? _T_23_mulres65_0 : PMDU1_bits_Pctrl_mulres65_0; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [65:0] _GEN_759 = PMDU1_io_in_ready ? _T_23_mulres33_0 : PMDU1_bits_Pctrl_mulres33_0; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [33:0] _GEN_760 = PMDU1_io_in_ready ? _T_23_mulres17_1 : PMDU1_bits_Pctrl_mulres17_1; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [33:0] _GEN_761 = PMDU1_io_in_ready ? _T_23_mulres17_0 : PMDU1_bits_Pctrl_mulres17_0; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [17:0] _GEN_762 = PMDU1_io_in_ready ? _T_23_mulres9_3 : PMDU1_bits_Pctrl_mulres9_3; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [17:0] _GEN_763 = PMDU1_io_in_ready ? _T_23_mulres9_2 : PMDU1_bits_Pctrl_mulres9_2; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [17:0] _GEN_764 = PMDU1_io_in_ready ? _T_23_mulres9_1 : PMDU1_bits_Pctrl_mulres9_1; // @[SIMDU.scala 508:19 539:34 543:32]
  wire [17:0] _GEN_765 = PMDU1_io_in_ready ? _T_23_mulres9_0 : PMDU1_bits_Pctrl_mulres9_0; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_766 = PMDU1_io_in_ready ? _T_23_isPMA_64ONLY : PMDU1_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_767 = PMDU1_io_in_ready ? _T_23_isMul_32_64ONLY : PMDU1_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_768 = PMDU1_io_in_ready ? _T_23_isQ63_64ONLY : PMDU1_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_769 = PMDU1_io_in_ready ? _T_23_isQ15_64ONLY : PMDU1_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_770 = PMDU1_io_in_ready ? _T_23_isC31 : PMDU1_bits_Pctrl_isC31; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_771 = PMDU1_io_in_ready ? _T_23_isQ15orQ31 : PMDU1_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_772 = PMDU1_io_in_ready ? _T_23_is1664 : PMDU1_bits_Pctrl_is1664; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_773 = PMDU1_io_in_ready ? _T_23_is3264 : PMDU1_bits_Pctrl_is3264; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_774 = PMDU1_io_in_ready ? _T_23_is832 : PMDU1_bits_Pctrl_is832; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_775 = PMDU1_io_in_ready ? _T_23_isS1664 : PMDU1_bits_Pctrl_isS1664; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_776 = PMDU1_io_in_ready ? _T_23_isS1632 : PMDU1_bits_Pctrl_isS1632; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_777 = PMDU1_io_in_ready ? _T_23_isMSW_3216 : PMDU1_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_778 = PMDU1_io_in_ready ? _T_23_isMSW_3232 : PMDU1_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_779 = PMDU1_io_in_ready ? _T_23_isMul_8 : PMDU1_bits_Pctrl_isMul_8; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_780 = PMDU1_io_in_ready ? _T_23_isMul_16 : PMDU1_bits_Pctrl_isMul_16; // @[SIMDU.scala 508:19 539:34 543:32]
  wire  _GEN_870 = PMDU1_io_in_ready & secondidx; // @[SIMDU.scala 472:24 539:34]
  wire  _GEN_871 = PMDU1_io_in_ready & firstidx; // @[SIMDU.scala 473:24 539:34]
  wire  _GEN_872 = PMDU0_io_in_ready; // @[SIMDU.scala 533:28 534:25]
  wire  _GEN_873 = PMDU0_io_in_ready | _GEN_2; // @[SIMDU.scala 533:28 535:24]
  wire  _GEN_874 = PMDU0_io_in_ready ? _GEN_9 : PMDU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [4:0] _GEN_875 = PMDU0_io_in_ready ? _GEN_11 : PMDU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [63:0] _GEN_878 = PMDU0_io_in_ready ? _GEN_17 : PMDU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [63:0] _GEN_879 = PMDU0_io_in_ready ? _GEN_19 : PMDU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [63:0] _GEN_880 = PMDU0_io_in_ready ? _GEN_21 : PMDU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [4:0] _GEN_888 = PMDU0_io_in_ready ? _GEN_37 : PMDU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 500:19 533:28 536:32]
  wire  _GEN_889 = PMDU0_io_in_ready ? _GEN_39 : PMDU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [6:0] _GEN_896 = PMDU0_io_in_ready ? _GEN_53 : PMDU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [63:0] _GEN_902 = PMDU0_io_in_ready ? _GEN_63 : PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [38:0] _GEN_938 = PMDU0_io_in_ready ? _GEN_135 : PMDU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 500:19 533:28 536:32]
  wire [129:0] _GEN_940 = PMDU0_io_in_ready ? _T_23_mulres65_0 : PMDU0_bits_Pctrl_mulres65_0; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [65:0] _GEN_941 = PMDU0_io_in_ready ? _T_23_mulres33_0 : PMDU0_bits_Pctrl_mulres33_0; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [33:0] _GEN_942 = PMDU0_io_in_ready ? _T_23_mulres17_1 : PMDU0_bits_Pctrl_mulres17_1; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [33:0] _GEN_943 = PMDU0_io_in_ready ? _T_23_mulres17_0 : PMDU0_bits_Pctrl_mulres17_0; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [17:0] _GEN_944 = PMDU0_io_in_ready ? _T_23_mulres9_3 : PMDU0_bits_Pctrl_mulres9_3; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [17:0] _GEN_945 = PMDU0_io_in_ready ? _T_23_mulres9_2 : PMDU0_bits_Pctrl_mulres9_2; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [17:0] _GEN_946 = PMDU0_io_in_ready ? _T_23_mulres9_1 : PMDU0_bits_Pctrl_mulres9_1; // @[SIMDU.scala 500:19 533:28 537:32]
  wire [17:0] _GEN_947 = PMDU0_io_in_ready ? _T_23_mulres9_0 : PMDU0_bits_Pctrl_mulres9_0; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_948 = PMDU0_io_in_ready ? _T_23_isPMA_64ONLY : PMDU0_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_949 = PMDU0_io_in_ready ? _T_23_isMul_32_64ONLY : PMDU0_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_950 = PMDU0_io_in_ready ? _T_23_isQ63_64ONLY : PMDU0_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_951 = PMDU0_io_in_ready ? _T_23_isQ15_64ONLY : PMDU0_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_952 = PMDU0_io_in_ready ? _T_23_isC31 : PMDU0_bits_Pctrl_isC31; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_953 = PMDU0_io_in_ready ? _T_23_isQ15orQ31 : PMDU0_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_954 = PMDU0_io_in_ready ? _T_23_is1664 : PMDU0_bits_Pctrl_is1664; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_955 = PMDU0_io_in_ready ? _T_23_is3264 : PMDU0_bits_Pctrl_is3264; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_956 = PMDU0_io_in_ready ? _T_23_is832 : PMDU0_bits_Pctrl_is832; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_957 = PMDU0_io_in_ready ? _T_23_isS1664 : PMDU0_bits_Pctrl_isS1664; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_958 = PMDU0_io_in_ready ? _T_23_isS1632 : PMDU0_bits_Pctrl_isS1632; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_959 = PMDU0_io_in_ready ? _T_23_isMSW_3216 : PMDU0_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_960 = PMDU0_io_in_ready ? _T_23_isMSW_3232 : PMDU0_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_961 = PMDU0_io_in_ready ? _T_23_isMul_8 : PMDU0_bits_Pctrl_isMul_8; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_962 = PMDU0_io_in_ready ? _T_23_isMul_16 : PMDU0_bits_Pctrl_isMul_16; // @[SIMDU.scala 500:19 533:28 537:32]
  wire  _GEN_1052 = PMDU0_io_in_ready ? secondidx : _GEN_870; // @[SIMDU.scala 533:28]
  wire  _GEN_1053 = PMDU0_io_in_ready ? firstidx : _GEN_871; // @[SIMDU.scala 533:28]
  wire  _GEN_1054 = PMDU0_io_in_ready ? 1'h0 : _GEN_690; // @[SIMDU.scala 533:28]
  wire  _GEN_1055 = PMDU0_io_in_ready ? _GEN_3 : _GEN_691; // @[SIMDU.scala 533:28]
  wire  _GEN_1056 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_InstFlag : _GEN_692; // @[SIMDU.scala 508:19 533:28]
  wire [4:0] _GEN_1057 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_InstNo : _GEN_693; // @[SIMDU.scala 508:19 533:28]
  wire [63:0] _GEN_1060 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_data_src3 : _GEN_696; // @[SIMDU.scala 508:19 533:28]
  wire [63:0] _GEN_1061 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_data_src2 : _GEN_697; // @[SIMDU.scala 508:19 533:28]
  wire [63:0] _GEN_1062 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_data_src1 : _GEN_698; // @[SIMDU.scala 508:19 533:28]
  wire [4:0] _GEN_1070 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_ctrl_rfDest : _GEN_706; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1071 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_ctrl_rfWen : _GEN_707; // @[SIMDU.scala 508:19 533:28]
  wire [6:0] _GEN_1078 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_ctrl_fuOpType : _GEN_714; // @[SIMDU.scala 508:19 533:28]
  wire [63:0] _GEN_1084 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id : _GEN_720; // @[SIMDU.scala 508:19 533:28]
  wire [38:0] _GEN_1120 = PMDU0_io_in_ready ? PMDU1_bits_DecodeIn_cf_pc : _GEN_756; // @[SIMDU.scala 508:19 533:28]
  wire [129:0] _GEN_1122 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres65_0 : _GEN_758; // @[SIMDU.scala 508:19 533:28]
  wire [65:0] _GEN_1123 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres33_0 : _GEN_759; // @[SIMDU.scala 508:19 533:28]
  wire [33:0] _GEN_1124 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres17_1 : _GEN_760; // @[SIMDU.scala 508:19 533:28]
  wire [33:0] _GEN_1125 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres17_0 : _GEN_761; // @[SIMDU.scala 508:19 533:28]
  wire [17:0] _GEN_1126 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres9_3 : _GEN_762; // @[SIMDU.scala 508:19 533:28]
  wire [17:0] _GEN_1127 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres9_2 : _GEN_763; // @[SIMDU.scala 508:19 533:28]
  wire [17:0] _GEN_1128 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres9_1 : _GEN_764; // @[SIMDU.scala 508:19 533:28]
  wire [17:0] _GEN_1129 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_mulres9_0 : _GEN_765; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1130 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isPMA_64ONLY : _GEN_766; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1131 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isMul_32_64ONLY : _GEN_767; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1132 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isQ63_64ONLY : _GEN_768; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1133 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isQ15_64ONLY : _GEN_769; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1134 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isC31 : _GEN_770; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1135 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isQ15orQ31 : _GEN_771; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1136 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_is1664 : _GEN_772; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1137 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_is3264 : _GEN_773; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1138 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_is832 : _GEN_774; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1139 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isS1664 : _GEN_775; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1140 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isS1632 : _GEN_776; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1141 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isMSW_3216 : _GEN_777; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1142 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isMSW_3232 : _GEN_778; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1143 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isMul_8 : _GEN_779; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1144 = PMDU0_io_in_ready ? PMDU1_bits_Pctrl_isMul_16 : _GEN_780; // @[SIMDU.scala 508:19 533:28]
  wire  _GEN_1234 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) & _GEN_872; // @[SIMDU.scala 532:139]
  wire  _GEN_1235 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_873 : _GEN_2; // @[SIMDU.scala 532:139]
  wire  _GEN_1236 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_874 : PMDU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 532:139 500:19]
  wire [4:0] _GEN_1237 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_875 : PMDU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 532:139 500:19]
  wire [63:0] _GEN_1240 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_878 : PMDU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 532:139 500:19]
  wire [63:0] _GEN_1241 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_879 : PMDU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 532:139 500:19]
  wire [63:0] _GEN_1242 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_880 : PMDU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 532:139 500:19]
  wire [4:0] _GEN_1250 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_888 : PMDU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1251 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_889 : PMDU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 532:139 500:19]
  wire [6:0] _GEN_1258 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_896 : PMDU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 532:139 500:19]
  wire [63:0] _GEN_1264 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_902 :
    PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 532:139 500:19]
  wire [38:0] _GEN_1300 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_938 : PMDU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 532:139 500:19]
  wire [129:0] _GEN_1302 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_940 : PMDU0_bits_Pctrl_mulres65_0; // @[SIMDU.scala 532:139 500:19]
  wire [65:0] _GEN_1303 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_941 : PMDU0_bits_Pctrl_mulres33_0; // @[SIMDU.scala 532:139 500:19]
  wire [33:0] _GEN_1304 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_942 : PMDU0_bits_Pctrl_mulres17_1; // @[SIMDU.scala 532:139 500:19]
  wire [33:0] _GEN_1305 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_943 : PMDU0_bits_Pctrl_mulres17_0; // @[SIMDU.scala 532:139 500:19]
  wire [17:0] _GEN_1306 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_944 : PMDU0_bits_Pctrl_mulres9_3; // @[SIMDU.scala 532:139 500:19]
  wire [17:0] _GEN_1307 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_945 : PMDU0_bits_Pctrl_mulres9_2; // @[SIMDU.scala 532:139 500:19]
  wire [17:0] _GEN_1308 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_946 : PMDU0_bits_Pctrl_mulres9_1; // @[SIMDU.scala 532:139 500:19]
  wire [17:0] _GEN_1309 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_947 : PMDU0_bits_Pctrl_mulres9_0; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1310 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_948 : PMDU0_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1311 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_949 : PMDU0_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1312 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_950 : PMDU0_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1313 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_951 : PMDU0_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1314 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_952 : PMDU0_bits_Pctrl_isC31; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1315 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_953 : PMDU0_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1316 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_954 : PMDU0_bits_Pctrl_is1664; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1317 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_955 : PMDU0_bits_Pctrl_is3264; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1318 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_956 : PMDU0_bits_Pctrl_is832; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1319 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_957 : PMDU0_bits_Pctrl_isS1664; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1320 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_958 : PMDU0_bits_Pctrl_isS1632; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1321 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_959 : PMDU0_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1322 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_960 : PMDU0_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1323 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_961 : PMDU0_bits_Pctrl_isMul_8; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1324 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_962 : PMDU0_bits_Pctrl_isMul_16; // @[SIMDU.scala 532:139 500:19]
  wire  _GEN_1414 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) & _GEN_1052; // @[SIMDU.scala 532:139 472:24]
  wire  _GEN_1415 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) & _GEN_1053; // @[SIMDU.scala 532:139 473:24]
  wire  _GEN_1416 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) & _GEN_1054; // @[SIMDU.scala 532:139]
  wire  _GEN_1417 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1055 : _GEN_3; // @[SIMDU.scala 532:139]
  wire  _GEN_1418 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1056 : PMDU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 532:139 508:19]
  wire [4:0] _GEN_1419 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1057 : PMDU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 532:139 508:19]
  wire [63:0] _GEN_1422 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1060 : PMDU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 532:139 508:19]
  wire [63:0] _GEN_1423 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1061 : PMDU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 532:139 508:19]
  wire [63:0] _GEN_1424 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1062 : PMDU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 532:139 508:19]
  wire [4:0] _GEN_1432 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1070 : PMDU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1433 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1071 : PMDU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 532:139 508:19]
  wire [6:0] _GEN_1440 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1078 : PMDU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 532:139 508:19]
  wire [63:0] _GEN_1446 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1084 :
    PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 532:139 508:19]
  wire [38:0] _GEN_1482 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1120 : PMDU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 532:139 508:19]
  wire [129:0] _GEN_1484 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1122 : PMDU1_bits_Pctrl_mulres65_0; // @[SIMDU.scala 532:139 508:19]
  wire [65:0] _GEN_1485 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1123 : PMDU1_bits_Pctrl_mulres33_0; // @[SIMDU.scala 532:139 508:19]
  wire [33:0] _GEN_1486 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1124 : PMDU1_bits_Pctrl_mulres17_1; // @[SIMDU.scala 532:139 508:19]
  wire [33:0] _GEN_1487 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1125 : PMDU1_bits_Pctrl_mulres17_0; // @[SIMDU.scala 532:139 508:19]
  wire [17:0] _GEN_1488 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1126 : PMDU1_bits_Pctrl_mulres9_3; // @[SIMDU.scala 532:139 508:19]
  wire [17:0] _GEN_1489 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1127 : PMDU1_bits_Pctrl_mulres9_2; // @[SIMDU.scala 532:139 508:19]
  wire [17:0] _GEN_1490 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1128 : PMDU1_bits_Pctrl_mulres9_1; // @[SIMDU.scala 532:139 508:19]
  wire [17:0] _GEN_1491 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1129 : PMDU1_bits_Pctrl_mulres9_0; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1492 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1130 : PMDU1_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1493 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1131 : PMDU1_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1494 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1132 : PMDU1_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1495 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1133 : PMDU1_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1496 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1134 : PMDU1_bits_Pctrl_isC31; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1497 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1135 : PMDU1_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1498 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1136 : PMDU1_bits_Pctrl_is1664; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1499 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1137 : PMDU1_bits_Pctrl_is3264; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1500 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1138 : PMDU1_bits_Pctrl_is832; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1501 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1139 : PMDU1_bits_Pctrl_isS1664; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1502 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1140 : PMDU1_bits_Pctrl_isS1632; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1503 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1141 : PMDU1_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1504 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1142 : PMDU1_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1505 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1143 : PMDU1_bits_Pctrl_isMul_8; // @[SIMDU.scala 532:139 508:19]
  wire  _GEN_1506 = _GEN_7 & (_GEN_5 == 5'h16 | _GEN_5 == 5'h1c) ? _GEN_1144 : PMDU1_bits_Pctrl_isMul_16; // @[SIMDU.scala 532:139 508:19]
  wire  match_operator_0 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) & _GEN_324; // @[SIMDU.scala 518:180]
  wire  _GEN_1597 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_325 : _GEN_0; // @[SIMDU.scala 518:180]
  wire  _GEN_1598 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_326 :
    PALU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 518:180 483:19]
  wire [4:0] _GEN_1599 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_327 :
    PALU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 518:180 483:19]
  wire [63:0] _GEN_1602 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_330 :
    PALU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 518:180 483:19]
  wire [63:0] _GEN_1603 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_331 :
    PALU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 518:180 483:19]
  wire [63:0] _GEN_1604 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_332 :
    PALU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 518:180 483:19]
  wire [4:0] _GEN_1612 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_340 :
    PALU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1613 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_341 :
    PALU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1618 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_346 :
    PALU0_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 518:180 483:19]
  wire [2:0] _GEN_1619 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_347 :
    PALU0_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 518:180 483:19]
  wire [6:0] _GEN_1620 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_348 :
    PALU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 518:180 483:19]
  wire [63:0] _GEN_1626 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_354 :
    PALU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 518:180 483:19]
  wire [38:0] _GEN_1662 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_390 :
    PALU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1687 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_415 :
    PALU0_bits_Pctrl_Arithmetic; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1688 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_416 :
    PALU0_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1689 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_417 : PALU0_bits_Pctrl_Round; // @[SIMDU.scala 518:180 483:19]
  wire [79:0] _GEN_1690 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_418 :
    PALU0_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 518:180 483:19]
  wire [63:0] _GEN_1691 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_419 :
    PALU0_bits_Pctrl_adderRes; // @[SIMDU.scala 518:180 483:19]
  wire [79:0] _GEN_1692 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_420 :
    PALU0_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1693 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_421 :
    PALU0_bits_Pctrl_LessThan; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1694 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_422 :
    PALU0_bits_Pctrl_LessEqual; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1695 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_423 :
    PALU0_bits_Pctrl_Translation; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1696 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_424 :
    PALU0_bits_Pctrl_Saturating; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1697 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_425 :
    PALU0_bits_Pctrl_SrcSigned; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1698 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_426 : PALU0_bits_Pctrl_isAdder
    ; // @[SIMDU.scala 518:180 483:19]
  wire [7:0] _GEN_1699 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_427 :
    PALU0_bits_Pctrl_isSub; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1700 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_428 : PALU0_bits_Pctrl_isPack; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1701 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_429 :
    PALU0_bits_Pctrl_isPacktt; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1702 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_430 :
    PALU0_bits_Pctrl_isPacktb; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1703 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_431 :
    PALU0_bits_Pctrl_isPackbt; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1704 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_432 :
    PALU0_bits_Pctrl_isPackbb; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1705 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_433 :
    PALU0_bits_Pctrl_isInsertb; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1706 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_434 : PALU0_bits_Pctrl_isCmix; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1707 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_435 :
    PALU0_bits_Pctrl_isBitrev; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1708 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_436 :
    PALU0_bits_Pctrl_isUnpack; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1709 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_437 : PALU0_bits_Pctrl_isSwap; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1710 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_438 :
    PALU0_bits_Pctrl_isSwap_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1711 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_439 :
    PALU0_bits_Pctrl_isSwap_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1712 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_440 : PALU0_bits_Pctrl_isCnt; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1713 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_441 :
    PALU0_bits_Pctrl_isCnt_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1714 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_442 : PALU0_bits_Pctrl_isCnt_8
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1715 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_443 :
    PALU0_bits_Pctrl_isCnt_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1716 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_444 : PALU0_bits_Pctrl_isSat; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1717 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_445 : PALU0_bits_Pctrl_isSat_W
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1718 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_446 :
    PALU0_bits_Pctrl_isSat_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1719 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_447 : PALU0_bits_Pctrl_isSat_8
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1720 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_448 :
    PALU0_bits_Pctrl_isSat_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1721 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_449 : PALU0_bits_Pctrl_isClip; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1722 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_450 :
    PALU0_bits_Pctrl_isclip_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1723 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_451 :
    PALU0_bits_Pctrl_isClip_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1724 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_452 :
    PALU0_bits_Pctrl_isClip_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1725 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_453 :
    PALU0_bits_Pctrl_isShifter; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1726 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_454 : PALU0_bits_Pctrl_isWext; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1727 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_455 : PALU0_bits_Pctrl_isFSRW; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1728 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_456 :
    PALU0_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1729 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_457 :
    PALU0_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1730 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_458 :
    PALU0_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1731 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_459 :
    PALU0_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1732 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_460 : PALU0_bits_Pctrl_isLR_32
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1733 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_461 : PALU0_bits_Pctrl_isLs_32
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1734 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_462 : PALU0_bits_Pctrl_isRs_32
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1735 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_463 : PALU0_bits_Pctrl_isLR_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1736 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_464 : PALU0_bits_Pctrl_isLs_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1737 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_465 : PALU0_bits_Pctrl_isRs_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1738 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_466 : PALU0_bits_Pctrl_isLR_16
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1739 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_467 : PALU0_bits_Pctrl_isLs_16
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1740 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_468 : PALU0_bits_Pctrl_isRs_16
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1741 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_469 : PALU0_bits_Pctrl_isPbs; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1742 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_470 :
    PALU0_bits_Pctrl_isMaxMin; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1743 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_471 :
    PALU0_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1744 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_472 :
    PALU0_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1745 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_473 :
    PALU0_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1746 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_474 :
    PALU0_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1747 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_475 :
    PALU0_bits_Pctrl_isCompare; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1748 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_476 :
    PALU0_bits_Pctrl_isComp_8; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1749 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_477 :
    PALU0_bits_Pctrl_isComp_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1751 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_479 :
    PALU0_bits_Pctrl_isStsa_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1752 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_480 :
    PALU0_bits_Pctrl_isStas_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1753 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_481 :
    PALU0_bits_Pctrl_isStsa_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1754 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_482 :
    PALU0_bits_Pctrl_isStas_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1756 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_484 :
    PALU0_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1757 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_485 :
    PALU0_bits_Pctrl_isCras_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1758 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_486 :
    PALU0_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1759 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_487 :
    PALU0_bits_Pctrl_isCras_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1760 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_488 :
    PALU0_bits_Pctrl_isSub_C31; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1761 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_489 :
    PALU0_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1762 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_490 :
    PALU0_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1763 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_491 : PALU0_bits_Pctrl_isSub_8
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1764 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_492 :
    PALU0_bits_Pctrl_isSub_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1765 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_493 :
    PALU0_bits_Pctrl_isSub_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1766 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_494 :
    PALU0_bits_Pctrl_isSub_64; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1768 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_496 : PALU0_bits_Pctrl_isAve; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1769 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_497 :
    PALU0_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1770 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_498 :
    PALU0_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1771 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_499 :
    PALU0_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1772 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_500 : PALU0_bits_Pctrl_isAdd_8
    ; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1773 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_501 :
    PALU0_bits_Pctrl_isAdd_16; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1774 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_502 :
    PALU0_bits_Pctrl_isAdd_32; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1775 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_503 :
    PALU0_bits_Pctrl_isAdd_64; // @[SIMDU.scala 518:180 483:19]
  wire  _GEN_1776 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_504 : _GEN_1414; // @[SIMDU.scala 518:180]
  wire  _GEN_1777 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_505 : _GEN_1415; // @[SIMDU.scala 518:180]
  wire  match_operator_1 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) & _GEN_506; // @[SIMDU.scala 518:180]
  wire  _GEN_1779 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_507 : _GEN_1; // @[SIMDU.scala 518:180]
  wire  _GEN_1780 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_508 :
    PALU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 518:180 491:19]
  wire [4:0] _GEN_1781 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_509 :
    PALU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 518:180 491:19]
  wire [63:0] _GEN_1784 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_512 :
    PALU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 518:180 491:19]
  wire [63:0] _GEN_1785 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_513 :
    PALU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 518:180 491:19]
  wire [63:0] _GEN_1786 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_514 :
    PALU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 518:180 491:19]
  wire [4:0] _GEN_1794 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_522 :
    PALU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1795 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_523 :
    PALU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1800 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_528 :
    PALU1_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 518:180 491:19]
  wire [2:0] _GEN_1801 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_529 :
    PALU1_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 518:180 491:19]
  wire [6:0] _GEN_1802 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_530 :
    PALU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 518:180 491:19]
  wire [63:0] _GEN_1808 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_536 :
    PALU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 518:180 491:19]
  wire [38:0] _GEN_1844 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_572 :
    PALU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1869 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_597 :
    PALU1_bits_Pctrl_Arithmetic; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1870 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_598 :
    PALU1_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1871 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_599 : PALU1_bits_Pctrl_Round; // @[SIMDU.scala 518:180 491:19]
  wire [79:0] _GEN_1872 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_600 :
    PALU1_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 518:180 491:19]
  wire [63:0] _GEN_1873 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_601 :
    PALU1_bits_Pctrl_adderRes; // @[SIMDU.scala 518:180 491:19]
  wire [79:0] _GEN_1874 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_602 :
    PALU1_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1875 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_603 :
    PALU1_bits_Pctrl_LessThan; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1876 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_604 :
    PALU1_bits_Pctrl_LessEqual; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1877 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_605 :
    PALU1_bits_Pctrl_Translation; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1878 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_606 :
    PALU1_bits_Pctrl_Saturating; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1879 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_607 :
    PALU1_bits_Pctrl_SrcSigned; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1880 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_608 : PALU1_bits_Pctrl_isAdder
    ; // @[SIMDU.scala 518:180 491:19]
  wire [7:0] _GEN_1881 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_609 :
    PALU1_bits_Pctrl_isSub; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1882 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_610 : PALU1_bits_Pctrl_isPack; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1883 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_611 :
    PALU1_bits_Pctrl_isPacktt; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1884 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_612 :
    PALU1_bits_Pctrl_isPacktb; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1885 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_613 :
    PALU1_bits_Pctrl_isPackbt; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1886 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_614 :
    PALU1_bits_Pctrl_isPackbb; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1887 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_615 :
    PALU1_bits_Pctrl_isInsertb; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1888 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_616 : PALU1_bits_Pctrl_isCmix; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1889 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_617 :
    PALU1_bits_Pctrl_isBitrev; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1890 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_618 :
    PALU1_bits_Pctrl_isUnpack; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1891 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_619 : PALU1_bits_Pctrl_isSwap; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1892 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_620 :
    PALU1_bits_Pctrl_isSwap_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1893 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_621 :
    PALU1_bits_Pctrl_isSwap_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1894 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_622 : PALU1_bits_Pctrl_isCnt; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1895 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_623 :
    PALU1_bits_Pctrl_isCnt_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1896 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_624 : PALU1_bits_Pctrl_isCnt_8
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1897 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_625 :
    PALU1_bits_Pctrl_isCnt_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1898 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_626 : PALU1_bits_Pctrl_isSat; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1899 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_627 : PALU1_bits_Pctrl_isSat_W
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1900 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_628 :
    PALU1_bits_Pctrl_isSat_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1901 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_629 : PALU1_bits_Pctrl_isSat_8
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1902 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_630 :
    PALU1_bits_Pctrl_isSat_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1903 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_631 : PALU1_bits_Pctrl_isClip; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1904 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_632 :
    PALU1_bits_Pctrl_isclip_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1905 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_633 :
    PALU1_bits_Pctrl_isClip_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1906 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_634 :
    PALU1_bits_Pctrl_isClip_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1907 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_635 :
    PALU1_bits_Pctrl_isShifter; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1908 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_636 : PALU1_bits_Pctrl_isWext; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1909 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_637 : PALU1_bits_Pctrl_isFSRW; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1910 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_638 :
    PALU1_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1911 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_639 :
    PALU1_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1912 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_640 :
    PALU1_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1913 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_641 :
    PALU1_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1914 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_642 : PALU1_bits_Pctrl_isLR_32
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1915 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_643 : PALU1_bits_Pctrl_isLs_32
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1916 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_644 : PALU1_bits_Pctrl_isRs_32
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1917 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_645 : PALU1_bits_Pctrl_isLR_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1918 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_646 : PALU1_bits_Pctrl_isLs_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1919 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_647 : PALU1_bits_Pctrl_isRs_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1920 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_648 : PALU1_bits_Pctrl_isLR_16
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1921 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_649 : PALU1_bits_Pctrl_isLs_16
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1922 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_650 : PALU1_bits_Pctrl_isRs_16
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1923 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_651 : PALU1_bits_Pctrl_isPbs; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1924 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_652 :
    PALU1_bits_Pctrl_isMaxMin; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1925 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_653 :
    PALU1_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1926 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_654 :
    PALU1_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1927 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_655 :
    PALU1_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1928 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_656 :
    PALU1_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1929 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_657 :
    PALU1_bits_Pctrl_isCompare; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1930 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_658 :
    PALU1_bits_Pctrl_isComp_8; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1931 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_659 :
    PALU1_bits_Pctrl_isComp_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1933 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_661 :
    PALU1_bits_Pctrl_isStsa_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1934 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_662 :
    PALU1_bits_Pctrl_isStas_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1935 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_663 :
    PALU1_bits_Pctrl_isStsa_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1936 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_664 :
    PALU1_bits_Pctrl_isStas_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1938 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_666 :
    PALU1_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1939 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_667 :
    PALU1_bits_Pctrl_isCras_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1940 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_668 :
    PALU1_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1941 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_669 :
    PALU1_bits_Pctrl_isCras_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1942 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_670 :
    PALU1_bits_Pctrl_isSub_C31; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1943 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_671 :
    PALU1_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1944 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_672 :
    PALU1_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1945 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_673 : PALU1_bits_Pctrl_isSub_8
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1946 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_674 :
    PALU1_bits_Pctrl_isSub_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1947 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_675 :
    PALU1_bits_Pctrl_isSub_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1948 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_676 :
    PALU1_bits_Pctrl_isSub_64; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1950 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_678 : PALU1_bits_Pctrl_isAve; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1951 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_679 :
    PALU1_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1952 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_680 :
    PALU1_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1953 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_681 :
    PALU1_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1954 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_682 : PALU1_bits_Pctrl_isAdd_8
    ; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1955 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_683 :
    PALU1_bits_Pctrl_isAdd_16; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1956 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_684 :
    PALU1_bits_Pctrl_isAdd_32; // @[SIMDU.scala 518:180 491:19]
  wire  _GEN_1957 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_685 :
    PALU1_bits_Pctrl_isAdd_64; // @[SIMDU.scala 518:180 491:19]
  wire  match_operator_2 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? 1'h0 : _GEN_1234; // @[SIMDU.scala 518:180]
  wire  _GEN_1959 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_2 : _GEN_1235; // @[SIMDU.scala 518:180]
  wire  _GEN_1960 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_InstFlag :
    _GEN_1236; // @[SIMDU.scala 518:180 500:19]
  wire [4:0] _GEN_1961 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_InstNo :
    _GEN_1237; // @[SIMDU.scala 518:180 500:19]
  wire [63:0] _GEN_1964 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_data_src3
     : _GEN_1240; // @[SIMDU.scala 518:180 500:19]
  wire [63:0] _GEN_1965 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_data_src2
     : _GEN_1241; // @[SIMDU.scala 518:180 500:19]
  wire [63:0] _GEN_1966 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_data_src1
     : _GEN_1242; // @[SIMDU.scala 518:180 500:19]
  wire [4:0] _GEN_1974 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ?
    PMDU0_bits_DecodeIn_ctrl_rfDest : _GEN_1250; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_1975 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_ctrl_rfWen :
    _GEN_1251; // @[SIMDU.scala 518:180 500:19]
  wire [6:0] _GEN_1982 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ?
    PMDU0_bits_DecodeIn_ctrl_fuOpType : _GEN_1258; // @[SIMDU.scala 518:180 500:19]
  wire [63:0] _GEN_1988 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ?
    PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id : _GEN_1264; // @[SIMDU.scala 518:180 500:19]
  wire [38:0] _GEN_2024 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_DecodeIn_cf_pc :
    _GEN_1300; // @[SIMDU.scala 518:180 500:19]
  wire [129:0] _GEN_2026 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres65_0
     : _GEN_1302; // @[SIMDU.scala 518:180 500:19]
  wire [65:0] _GEN_2027 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres33_0
     : _GEN_1303; // @[SIMDU.scala 518:180 500:19]
  wire [33:0] _GEN_2028 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres17_1
     : _GEN_1304; // @[SIMDU.scala 518:180 500:19]
  wire [33:0] _GEN_2029 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres17_0
     : _GEN_1305; // @[SIMDU.scala 518:180 500:19]
  wire [17:0] _GEN_2030 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres9_3 :
    _GEN_1306; // @[SIMDU.scala 518:180 500:19]
  wire [17:0] _GEN_2031 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres9_2 :
    _GEN_1307; // @[SIMDU.scala 518:180 500:19]
  wire [17:0] _GEN_2032 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres9_1 :
    _GEN_1308; // @[SIMDU.scala 518:180 500:19]
  wire [17:0] _GEN_2033 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_mulres9_0 :
    _GEN_1309; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2034 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isPMA_64ONLY :
    _GEN_1310; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2035 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isMul_32_64ONLY :
    _GEN_1311; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2036 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isQ63_64ONLY :
    _GEN_1312; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2037 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isQ15_64ONLY :
    _GEN_1313; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2038 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isC31 : _GEN_1314; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2039 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isQ15orQ31 :
    _GEN_1315; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2040 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_is1664 : _GEN_1316
    ; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2041 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_is3264 : _GEN_1317
    ; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2042 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_is832 : _GEN_1318; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2043 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isS1664 :
    _GEN_1319; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2044 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isS1632 :
    _GEN_1320; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2045 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isMSW_3216 :
    _GEN_1321; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2046 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isMSW_3232 :
    _GEN_1322; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2047 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isMul_8 :
    _GEN_1323; // @[SIMDU.scala 518:180 500:19]
  wire  _GEN_2048 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU0_bits_Pctrl_isMul_16 :
    _GEN_1324; // @[SIMDU.scala 518:180 500:19]
  wire  match_operator_3 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? 1'h0 : _GEN_1416; // @[SIMDU.scala 518:180]
  wire  _GEN_2139 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? _GEN_3 : _GEN_1417; // @[SIMDU.scala 518:180]
  wire  _GEN_2140 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_InstFlag :
    _GEN_1418; // @[SIMDU.scala 518:180 508:19]
  wire [4:0] _GEN_2141 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_InstNo :
    _GEN_1419; // @[SIMDU.scala 518:180 508:19]
  wire [63:0] _GEN_2144 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_data_src3
     : _GEN_1422; // @[SIMDU.scala 518:180 508:19]
  wire [63:0] _GEN_2145 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_data_src2
     : _GEN_1423; // @[SIMDU.scala 518:180 508:19]
  wire [63:0] _GEN_2146 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_data_src1
     : _GEN_1424; // @[SIMDU.scala 518:180 508:19]
  wire [4:0] _GEN_2154 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ?
    PMDU1_bits_DecodeIn_ctrl_rfDest : _GEN_1432; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2155 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_ctrl_rfWen :
    _GEN_1433; // @[SIMDU.scala 518:180 508:19]
  wire [6:0] _GEN_2162 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ?
    PMDU1_bits_DecodeIn_ctrl_fuOpType : _GEN_1440; // @[SIMDU.scala 518:180 508:19]
  wire [63:0] _GEN_2168 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ?
    PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id : _GEN_1446; // @[SIMDU.scala 518:180 508:19]
  wire [38:0] _GEN_2204 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_DecodeIn_cf_pc :
    _GEN_1482; // @[SIMDU.scala 518:180 508:19]
  wire [129:0] _GEN_2206 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres65_0
     : _GEN_1484; // @[SIMDU.scala 518:180 508:19]
  wire [65:0] _GEN_2207 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres33_0
     : _GEN_1485; // @[SIMDU.scala 518:180 508:19]
  wire [33:0] _GEN_2208 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres17_1
     : _GEN_1486; // @[SIMDU.scala 518:180 508:19]
  wire [33:0] _GEN_2209 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres17_0
     : _GEN_1487; // @[SIMDU.scala 518:180 508:19]
  wire [17:0] _GEN_2210 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres9_3 :
    _GEN_1488; // @[SIMDU.scala 518:180 508:19]
  wire [17:0] _GEN_2211 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres9_2 :
    _GEN_1489; // @[SIMDU.scala 518:180 508:19]
  wire [17:0] _GEN_2212 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres9_1 :
    _GEN_1490; // @[SIMDU.scala 518:180 508:19]
  wire [17:0] _GEN_2213 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_mulres9_0 :
    _GEN_1491; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2214 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isPMA_64ONLY :
    _GEN_1492; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2215 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isMul_32_64ONLY :
    _GEN_1493; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2216 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isQ63_64ONLY :
    _GEN_1494; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2217 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isQ15_64ONLY :
    _GEN_1495; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2218 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isC31 : _GEN_1496; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2219 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isQ15orQ31 :
    _GEN_1497; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2220 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_is1664 : _GEN_1498
    ; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2221 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_is3264 : _GEN_1499
    ; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2222 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_is832 : _GEN_1500; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2223 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isS1664 :
    _GEN_1501; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2224 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isS1632 :
    _GEN_1502; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2225 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isMSW_3216 :
    _GEN_1503; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2226 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isMSW_3232 :
    _GEN_1504; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2227 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isMul_8 :
    _GEN_1505; // @[SIMDU.scala 518:180 508:19]
  wire  _GEN_2228 = _GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15) ? PMDU1_bits_Pctrl_isMul_16 :
    _GEN_1506; // @[SIMDU.scala 518:180 508:19]
  wire [4:0] _GEN_2319 = secondidx ? io_DecodeIn_1_cf_instrType : io_DecodeIn_0_cf_instrType; // @[SIMDU.scala 547:{71,71}]
  wire  _GEN_2321 = secondidx ? io_in_1_valid : io_in_0_valid; // @[SIMDU.scala 547:{31,31}]
  wire  _GEN_2323 = secondidx ? io_DecodeIn_1_InstFlag : io_DecodeIn_0_InstFlag; // @[SIMDU.scala 550:{32,32}]
  wire [4:0] _GEN_2325 = secondidx ? io_DecodeIn_1_InstNo : io_DecodeIn_0_InstNo; // @[SIMDU.scala 550:{32,32}]
  wire [63:0] _GEN_2331 = secondidx ? io_DecodeIn_1_data_src3 : io_DecodeIn_0_data_src3; // @[SIMDU.scala 550:{32,32}]
  wire [63:0] _GEN_2333 = secondidx ? io_DecodeIn_1_data_src2 : io_DecodeIn_0_data_src2; // @[SIMDU.scala 550:{32,32}]
  wire [63:0] _GEN_2335 = secondidx ? io_DecodeIn_1_data_src1 : io_DecodeIn_0_data_src1; // @[SIMDU.scala 550:{32,32}]
  wire [4:0] _GEN_2351 = secondidx ? io_DecodeIn_1_ctrl_rfDest : io_DecodeIn_0_ctrl_rfDest; // @[SIMDU.scala 550:{32,32}]
  wire  _GEN_2353 = secondidx ? io_DecodeIn_1_ctrl_rfWen : io_DecodeIn_0_ctrl_rfWen; // @[SIMDU.scala 550:{32,32}]
  wire  _GEN_2363 = secondidx ? io_DecodeIn_1_ctrl_func24 : io_DecodeIn_0_ctrl_func24; // @[SIMDU.scala 550:{32,32}]
  wire [2:0] _GEN_2365 = secondidx ? io_DecodeIn_1_ctrl_funct3 : io_DecodeIn_0_ctrl_funct3; // @[SIMDU.scala 550:{32,32}]
  wire [6:0] _GEN_2367 = secondidx ? io_DecodeIn_1_ctrl_fuOpType : io_DecodeIn_0_ctrl_fuOpType; // @[SIMDU.scala 550:{32,32}]
  wire [63:0] _GEN_2377 = secondidx ? io_DecodeIn_1_cf_runahead_checkpoint_id : io_DecodeIn_0_cf_runahead_checkpoint_id; // @[SIMDU.scala 550:{32,32}]
  wire [38:0] _GEN_2449 = secondidx ? io_DecodeIn_1_cf_pc : io_DecodeIn_0_cf_pc; // @[SIMDU.scala 550:{32,32}]
  wire  _T_42 = ~secondidx; // @[SIMDU.scala 551:49]
  wire  _T_43_isAdd_64 = ~secondidx ? PIDU0_io_Pctrl_isAdd_64 : PIDU1_io_Pctrl_isAdd_64; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdd_32 = ~secondidx ? PIDU0_io_Pctrl_isAdd_32 : PIDU1_io_Pctrl_isAdd_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdd_16 = ~secondidx ? PIDU0_io_Pctrl_isAdd_16 : PIDU1_io_Pctrl_isAdd_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdd_8 = ~secondidx ? PIDU0_io_Pctrl_isAdd_8 : PIDU1_io_Pctrl_isAdd_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdd_Q15 = ~secondidx ? PIDU0_io_Pctrl_isAdd_Q15 : PIDU1_io_Pctrl_isAdd_Q15; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdd_Q31 = ~secondidx ? PIDU0_io_Pctrl_isAdd_Q31 : PIDU1_io_Pctrl_isAdd_Q31; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdd_C31 = ~secondidx ? PIDU0_io_Pctrl_isAdd_C31 : PIDU1_io_Pctrl_isAdd_C31; // @[SIMDU.scala 551:38]
  wire  _T_43_isAve = ~secondidx ? PIDU0_io_Pctrl_isAve : PIDU1_io_Pctrl_isAve; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_64 = ~secondidx ? PIDU0_io_Pctrl_isSub_64 : PIDU1_io_Pctrl_isSub_64; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_32 = ~secondidx ? PIDU0_io_Pctrl_isSub_32 : PIDU1_io_Pctrl_isSub_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_16 = ~secondidx ? PIDU0_io_Pctrl_isSub_16 : PIDU1_io_Pctrl_isSub_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_8 = ~secondidx ? PIDU0_io_Pctrl_isSub_8 : PIDU1_io_Pctrl_isSub_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_Q15 = ~secondidx ? PIDU0_io_Pctrl_isSub_Q15 : PIDU1_io_Pctrl_isSub_Q15; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_Q31 = ~secondidx ? PIDU0_io_Pctrl_isSub_Q31 : PIDU1_io_Pctrl_isSub_Q31; // @[SIMDU.scala 551:38]
  wire  _T_43_isSub_C31 = ~secondidx ? PIDU0_io_Pctrl_isSub_C31 : PIDU1_io_Pctrl_isSub_C31; // @[SIMDU.scala 551:38]
  wire  _T_43_isCras_16 = ~secondidx ? PIDU0_io_Pctrl_isCras_16 : PIDU1_io_Pctrl_isCras_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isCrsa_16 = ~secondidx ? PIDU0_io_Pctrl_isCrsa_16 : PIDU1_io_Pctrl_isCrsa_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isCras_32 = ~secondidx ? PIDU0_io_Pctrl_isCras_32 : PIDU1_io_Pctrl_isCras_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isCrsa_32 = ~secondidx ? PIDU0_io_Pctrl_isCrsa_32 : PIDU1_io_Pctrl_isCrsa_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isStas_16 = ~secondidx ? PIDU0_io_Pctrl_isStas_16 : PIDU1_io_Pctrl_isStas_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isStsa_16 = ~secondidx ? PIDU0_io_Pctrl_isStsa_16 : PIDU1_io_Pctrl_isStsa_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isStas_32 = ~secondidx ? PIDU0_io_Pctrl_isStas_32 : PIDU1_io_Pctrl_isStas_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isStsa_32 = ~secondidx ? PIDU0_io_Pctrl_isStsa_32 : PIDU1_io_Pctrl_isStsa_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isComp_16 = ~secondidx ? PIDU0_io_Pctrl_isComp_16 : PIDU1_io_Pctrl_isComp_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isComp_8 = ~secondidx ? PIDU0_io_Pctrl_isComp_8 : PIDU1_io_Pctrl_isComp_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isCompare = ~secondidx ? PIDU0_io_Pctrl_isCompare : PIDU1_io_Pctrl_isCompare; // @[SIMDU.scala 551:38]
  wire  _T_43_isMaxMin_16 = ~secondidx ? PIDU0_io_Pctrl_isMaxMin_16 : PIDU1_io_Pctrl_isMaxMin_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isMaxMin_8 = ~secondidx ? PIDU0_io_Pctrl_isMaxMin_8 : PIDU1_io_Pctrl_isMaxMin_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isMaxMin_XLEN = ~secondidx ? PIDU0_io_Pctrl_isMaxMin_XLEN : PIDU1_io_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 551:38]
  wire  _T_43_isMaxMin_32 = ~secondidx ? PIDU0_io_Pctrl_isMaxMin_32 : PIDU1_io_Pctrl_isMaxMin_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isMaxMin = ~secondidx ? PIDU0_io_Pctrl_isMaxMin : PIDU1_io_Pctrl_isMaxMin; // @[SIMDU.scala 551:38]
  wire  _T_43_isPbs = ~secondidx ? PIDU0_io_Pctrl_isPbs : PIDU1_io_Pctrl_isPbs; // @[SIMDU.scala 551:38]
  wire  _T_43_isRs_16 = ~secondidx ? PIDU0_io_Pctrl_isRs_16 : PIDU1_io_Pctrl_isRs_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isLs_16 = ~secondidx ? PIDU0_io_Pctrl_isLs_16 : PIDU1_io_Pctrl_isLs_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isLR_16 = ~secondidx ? PIDU0_io_Pctrl_isLR_16 : PIDU1_io_Pctrl_isLR_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isRs_8 = ~secondidx ? PIDU0_io_Pctrl_isRs_8 : PIDU1_io_Pctrl_isRs_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isLs_8 = ~secondidx ? PIDU0_io_Pctrl_isLs_8 : PIDU1_io_Pctrl_isLs_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isLR_8 = ~secondidx ? PIDU0_io_Pctrl_isLR_8 : PIDU1_io_Pctrl_isLR_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isRs_32 = ~secondidx ? PIDU0_io_Pctrl_isRs_32 : PIDU1_io_Pctrl_isRs_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isLs_32 = ~secondidx ? PIDU0_io_Pctrl_isLs_32 : PIDU1_io_Pctrl_isLs_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isLR_32 = ~secondidx ? PIDU0_io_Pctrl_isLR_32 : PIDU1_io_Pctrl_isLR_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isLR_Q31 = ~secondidx ? PIDU0_io_Pctrl_isLR_Q31 : PIDU1_io_Pctrl_isLR_Q31; // @[SIMDU.scala 551:38]
  wire  _T_43_isLs_Q31 = ~secondidx ? PIDU0_io_Pctrl_isLs_Q31 : PIDU1_io_Pctrl_isLs_Q31; // @[SIMDU.scala 551:38]
  wire  _T_43_isRs_XLEN = ~secondidx ? PIDU0_io_Pctrl_isRs_XLEN : PIDU1_io_Pctrl_isRs_XLEN; // @[SIMDU.scala 551:38]
  wire  _T_43_isSRAIWU = ~secondidx ? PIDU0_io_Pctrl_isSRAIWU : PIDU1_io_Pctrl_isSRAIWU; // @[SIMDU.scala 551:38]
  wire  _T_43_isFSRW = ~secondidx ? PIDU0_io_Pctrl_isFSRW : PIDU1_io_Pctrl_isFSRW; // @[SIMDU.scala 551:38]
  wire  _T_43_isWext = ~secondidx ? PIDU0_io_Pctrl_isWext : PIDU1_io_Pctrl_isWext; // @[SIMDU.scala 551:38]
  wire  _T_43_isShifter = ~secondidx ? PIDU0_io_Pctrl_isShifter : PIDU1_io_Pctrl_isShifter; // @[SIMDU.scala 551:38]
  wire  _T_43_isClip_16 = ~secondidx ? PIDU0_io_Pctrl_isClip_16 : PIDU1_io_Pctrl_isClip_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isClip_8 = ~secondidx ? PIDU0_io_Pctrl_isClip_8 : PIDU1_io_Pctrl_isClip_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isclip_32 = ~secondidx ? PIDU0_io_Pctrl_isclip_32 : PIDU1_io_Pctrl_isclip_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isClip = ~secondidx ? PIDU0_io_Pctrl_isClip : PIDU1_io_Pctrl_isClip; // @[SIMDU.scala 551:38]
  wire  _T_43_isSat_16 = ~secondidx ? PIDU0_io_Pctrl_isSat_16 : PIDU1_io_Pctrl_isSat_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isSat_8 = ~secondidx ? PIDU0_io_Pctrl_isSat_8 : PIDU1_io_Pctrl_isSat_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isSat_32 = ~secondidx ? PIDU0_io_Pctrl_isSat_32 : PIDU1_io_Pctrl_isSat_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isSat_W = ~secondidx ? PIDU0_io_Pctrl_isSat_W : PIDU1_io_Pctrl_isSat_W; // @[SIMDU.scala 551:38]
  wire  _T_43_isSat = ~secondidx ? PIDU0_io_Pctrl_isSat : PIDU1_io_Pctrl_isSat; // @[SIMDU.scala 551:38]
  wire  _T_43_isCnt_16 = ~secondidx ? PIDU0_io_Pctrl_isCnt_16 : PIDU1_io_Pctrl_isCnt_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isCnt_8 = ~secondidx ? PIDU0_io_Pctrl_isCnt_8 : PIDU1_io_Pctrl_isCnt_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isCnt_32 = ~secondidx ? PIDU0_io_Pctrl_isCnt_32 : PIDU1_io_Pctrl_isCnt_32; // @[SIMDU.scala 551:38]
  wire  _T_43_isCnt = ~secondidx ? PIDU0_io_Pctrl_isCnt : PIDU1_io_Pctrl_isCnt; // @[SIMDU.scala 551:38]
  wire  _T_43_isSwap_16 = ~secondidx ? PIDU0_io_Pctrl_isSwap_16 : PIDU1_io_Pctrl_isSwap_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isSwap_8 = ~secondidx ? PIDU0_io_Pctrl_isSwap_8 : PIDU1_io_Pctrl_isSwap_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isSwap = ~secondidx ? PIDU0_io_Pctrl_isSwap : PIDU1_io_Pctrl_isSwap; // @[SIMDU.scala 551:38]
  wire  _T_43_isUnpack = ~secondidx ? PIDU0_io_Pctrl_isUnpack : PIDU1_io_Pctrl_isUnpack; // @[SIMDU.scala 551:38]
  wire  _T_43_isBitrev = ~secondidx ? PIDU0_io_Pctrl_isBitrev : PIDU1_io_Pctrl_isBitrev; // @[SIMDU.scala 551:38]
  wire  _T_43_isCmix = ~secondidx ? PIDU0_io_Pctrl_isCmix : PIDU1_io_Pctrl_isCmix; // @[SIMDU.scala 551:38]
  wire  _T_43_isInsertb = ~secondidx ? PIDU0_io_Pctrl_isInsertb : PIDU1_io_Pctrl_isInsertb; // @[SIMDU.scala 551:38]
  wire  _T_43_isPackbb = ~secondidx ? PIDU0_io_Pctrl_isPackbb : PIDU1_io_Pctrl_isPackbb; // @[SIMDU.scala 551:38]
  wire  _T_43_isPackbt = ~secondidx ? PIDU0_io_Pctrl_isPackbt : PIDU1_io_Pctrl_isPackbt; // @[SIMDU.scala 551:38]
  wire  _T_43_isPacktb = ~secondidx ? PIDU0_io_Pctrl_isPacktb : PIDU1_io_Pctrl_isPacktb; // @[SIMDU.scala 551:38]
  wire  _T_43_isPacktt = ~secondidx ? PIDU0_io_Pctrl_isPacktt : PIDU1_io_Pctrl_isPacktt; // @[SIMDU.scala 551:38]
  wire  _T_43_isPack = ~secondidx ? PIDU0_io_Pctrl_isPack : PIDU1_io_Pctrl_isPack; // @[SIMDU.scala 551:38]
  wire [7:0] _T_43_isSub = ~secondidx ? PIDU0_io_Pctrl_isSub : PIDU1_io_Pctrl_isSub; // @[SIMDU.scala 551:38]
  wire  _T_43_isAdder = ~secondidx ? PIDU0_io_Pctrl_isAdder : PIDU1_io_Pctrl_isAdder; // @[SIMDU.scala 551:38]
  wire  _T_43_SrcSigned = ~secondidx ? PIDU0_io_Pctrl_SrcSigned : PIDU1_io_Pctrl_SrcSigned; // @[SIMDU.scala 551:38]
  wire  _T_43_Saturating = ~secondidx ? PIDU0_io_Pctrl_Saturating : PIDU1_io_Pctrl_Saturating; // @[SIMDU.scala 551:38]
  wire  _T_43_Translation = ~secondidx ? PIDU0_io_Pctrl_Translation : PIDU1_io_Pctrl_Translation; // @[SIMDU.scala 551:38]
  wire  _T_43_LessEqual = ~secondidx ? PIDU0_io_Pctrl_LessEqual : PIDU1_io_Pctrl_LessEqual; // @[SIMDU.scala 551:38]
  wire  _T_43_LessThan = ~secondidx ? PIDU0_io_Pctrl_LessThan : PIDU1_io_Pctrl_LessThan; // @[SIMDU.scala 551:38]
  wire [79:0] _T_43_adderRes_ori = ~secondidx ? PIDU0_io_Pctrl_adderRes_ori : PIDU1_io_Pctrl_adderRes_ori; // @[SIMDU.scala 551:38]
  wire [63:0] _T_43_adderRes = ~secondidx ? PIDU0_io_Pctrl_adderRes : PIDU1_io_Pctrl_adderRes; // @[SIMDU.scala 551:38]
  wire [79:0] _T_43_adderRes_ori_drophighestbit = ~secondidx ? PIDU0_io_Pctrl_adderRes_ori_drophighestbit :
    PIDU1_io_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 551:38]
  wire  _T_43_Round = ~secondidx ? PIDU0_io_Pctrl_Round : PIDU1_io_Pctrl_Round; // @[SIMDU.scala 551:38]
  wire  _T_43_ShiftSigned = ~secondidx ? PIDU0_io_Pctrl_ShiftSigned : PIDU1_io_Pctrl_ShiftSigned; // @[SIMDU.scala 551:38]
  wire  _T_43_Arithmetic = ~secondidx ? PIDU0_io_Pctrl_Arithmetic : PIDU1_io_Pctrl_Arithmetic; // @[SIMDU.scala 551:38]
  wire  _T_43_isMul_16 = ~secondidx ? PIDU0_io_Pctrl_isMul_16 : PIDU1_io_Pctrl_isMul_16; // @[SIMDU.scala 551:38]
  wire  _T_43_isMul_8 = ~secondidx ? PIDU0_io_Pctrl_isMul_8 : PIDU1_io_Pctrl_isMul_8; // @[SIMDU.scala 551:38]
  wire  _T_43_isMSW_3232 = ~secondidx ? PIDU0_io_Pctrl_isMSW_3232 : PIDU1_io_Pctrl_isMSW_3232; // @[SIMDU.scala 551:38]
  wire  _T_43_isMSW_3216 = ~secondidx ? PIDU0_io_Pctrl_isMSW_3216 : PIDU1_io_Pctrl_isMSW_3216; // @[SIMDU.scala 551:38]
  wire  _T_43_isS1632 = ~secondidx ? PIDU0_io_Pctrl_isS1632 : PIDU1_io_Pctrl_isS1632; // @[SIMDU.scala 551:38]
  wire  _T_43_isS1664 = ~secondidx ? PIDU0_io_Pctrl_isS1664 : PIDU1_io_Pctrl_isS1664; // @[SIMDU.scala 551:38]
  wire  _T_43_is832 = ~secondidx ? PIDU0_io_Pctrl_is832 : PIDU1_io_Pctrl_is832; // @[SIMDU.scala 551:38]
  wire  _T_43_is3264 = ~secondidx ? PIDU0_io_Pctrl_is3264 : PIDU1_io_Pctrl_is3264; // @[SIMDU.scala 551:38]
  wire  _T_43_is1664 = ~secondidx ? PIDU0_io_Pctrl_is1664 : PIDU1_io_Pctrl_is1664; // @[SIMDU.scala 551:38]
  wire  _T_43_isQ15orQ31 = ~secondidx ? PIDU0_io_Pctrl_isQ15orQ31 : PIDU1_io_Pctrl_isQ15orQ31; // @[SIMDU.scala 551:38]
  wire  _T_43_isC31 = ~secondidx ? PIDU0_io_Pctrl_isC31 : PIDU1_io_Pctrl_isC31; // @[SIMDU.scala 551:38]
  wire  _T_43_isQ15_64ONLY = ~secondidx ? PIDU0_io_Pctrl_isQ15_64ONLY : PIDU1_io_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 551:38]
  wire  _T_43_isQ63_64ONLY = ~secondidx ? PIDU0_io_Pctrl_isQ63_64ONLY : PIDU1_io_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 551:38]
  wire  _T_43_isMul_32_64ONLY = ~secondidx ? PIDU0_io_Pctrl_isMul_32_64ONLY : PIDU1_io_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 551:38]
  wire  _T_43_isPMA_64ONLY = ~secondidx ? PIDU0_io_Pctrl_isPMA_64ONLY : PIDU1_io_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 551:38]
  wire [17:0] _T_43_mulres9_0 = ~secondidx ? PIDU0_io_Pctrl_mulres9_0 : PIDU1_io_Pctrl_mulres9_0; // @[SIMDU.scala 551:38]
  wire [17:0] _T_43_mulres9_1 = ~secondidx ? PIDU0_io_Pctrl_mulres9_1 : PIDU1_io_Pctrl_mulres9_1; // @[SIMDU.scala 551:38]
  wire [17:0] _T_43_mulres9_2 = ~secondidx ? PIDU0_io_Pctrl_mulres9_2 : PIDU1_io_Pctrl_mulres9_2; // @[SIMDU.scala 551:38]
  wire [17:0] _T_43_mulres9_3 = ~secondidx ? PIDU0_io_Pctrl_mulres9_3 : PIDU1_io_Pctrl_mulres9_3; // @[SIMDU.scala 551:38]
  wire [33:0] _T_43_mulres17_0 = ~secondidx ? PIDU0_io_Pctrl_mulres17_0 : PIDU1_io_Pctrl_mulres17_0; // @[SIMDU.scala 551:38]
  wire [33:0] _T_43_mulres17_1 = ~secondidx ? PIDU0_io_Pctrl_mulres17_1 : PIDU1_io_Pctrl_mulres17_1; // @[SIMDU.scala 551:38]
  wire [65:0] _T_43_mulres33_0 = ~secondidx ? PIDU0_io_Pctrl_mulres33_0 : PIDU1_io_Pctrl_mulres33_0; // @[SIMDU.scala 551:38]
  wire [129:0] _T_43_mulres65_0 = ~secondidx ? PIDU0_io_Pctrl_mulres65_0 : PIDU1_io_Pctrl_mulres65_0; // @[SIMDU.scala 551:38]
  wire  _GEN_2452 = _T_42 | _GEN_1776; // @[SIMDU.scala 552:{36,36}]
  wire  _GEN_2453 = secondidx | _GEN_1777; // @[SIMDU.scala 552:{36,36}]
  wire  _GEN_2456 = PALU1_io_in_ready & ~match_operator_1 | _GEN_1779; // @[SIMDU.scala 553:56 554:24]
  wire  _GEN_2635 = PALU1_io_in_ready & ~match_operator_1 ? _GEN_2452 : _GEN_1776; // @[SIMDU.scala 553:56]
  wire  _GEN_2636 = PALU1_io_in_ready & ~match_operator_1 ? _GEN_2453 : _GEN_1777; // @[SIMDU.scala 553:56]
  wire  _GEN_2637 = PALU0_io_in_ready & ~match_operator_0 | _GEN_1597; // @[SIMDU.scala 548:50 549:24]
  wire  _GEN_2816 = PALU0_io_in_ready & ~match_operator_0 ? _GEN_2452 : _GEN_2635; // @[SIMDU.scala 548:50]
  wire  _GEN_2817 = PALU0_io_in_ready & ~match_operator_0 ? _GEN_2453 : _GEN_2636; // @[SIMDU.scala 548:50]
  wire  _GEN_3001 = PMDU1_io_in_ready & ~match_operator_3 | _GEN_2139; // @[SIMDU.scala 565:56 566:24]
  wire  _GEN_3002 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2323 : _GEN_2140; // @[SIMDU.scala 565:56 567:32]
  wire [4:0] _GEN_3003 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2325 : _GEN_2141; // @[SIMDU.scala 565:56 567:32]
  wire [63:0] _GEN_3006 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2331 : _GEN_2144; // @[SIMDU.scala 565:56 567:32]
  wire [63:0] _GEN_3007 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2333 : _GEN_2145; // @[SIMDU.scala 565:56 567:32]
  wire [63:0] _GEN_3008 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2335 : _GEN_2146; // @[SIMDU.scala 565:56 567:32]
  wire [4:0] _GEN_3016 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2351 : _GEN_2154; // @[SIMDU.scala 565:56 567:32]
  wire  _GEN_3017 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2353 : _GEN_2155; // @[SIMDU.scala 565:56 567:32]
  wire [6:0] _GEN_3024 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2367 : _GEN_2162; // @[SIMDU.scala 565:56 567:32]
  wire [63:0] _GEN_3030 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2377 : _GEN_2168; // @[SIMDU.scala 565:56 567:32]
  wire [38:0] _GEN_3066 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2449 : _GEN_2204; // @[SIMDU.scala 565:56 567:32]
  wire [129:0] _GEN_3068 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres65_0 : _GEN_2206; // @[SIMDU.scala 565:56 568:32]
  wire [65:0] _GEN_3069 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres33_0 : _GEN_2207; // @[SIMDU.scala 565:56 568:32]
  wire [33:0] _GEN_3070 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres17_1 : _GEN_2208; // @[SIMDU.scala 565:56 568:32]
  wire [33:0] _GEN_3071 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres17_0 : _GEN_2209; // @[SIMDU.scala 565:56 568:32]
  wire [17:0] _GEN_3072 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres9_3 : _GEN_2210; // @[SIMDU.scala 565:56 568:32]
  wire [17:0] _GEN_3073 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres9_2 : _GEN_2211; // @[SIMDU.scala 565:56 568:32]
  wire [17:0] _GEN_3074 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres9_1 : _GEN_2212; // @[SIMDU.scala 565:56 568:32]
  wire [17:0] _GEN_3075 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_mulres9_0 : _GEN_2213; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3076 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isPMA_64ONLY : _GEN_2214; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3077 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isMul_32_64ONLY : _GEN_2215; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3078 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isQ63_64ONLY : _GEN_2216; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3079 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isQ15_64ONLY : _GEN_2217; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3080 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isC31 : _GEN_2218; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3081 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isQ15orQ31 : _GEN_2219; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3082 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_is1664 : _GEN_2220; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3083 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_is3264 : _GEN_2221; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3084 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_is832 : _GEN_2222; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3085 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isS1664 : _GEN_2223; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3086 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isS1632 : _GEN_2224; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3087 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isMSW_3216 : _GEN_2225; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3088 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isMSW_3232 : _GEN_2226; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3089 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isMul_8 : _GEN_2227; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3090 = PMDU1_io_in_ready & ~match_operator_3 ? _T_43_isMul_16 : _GEN_2228; // @[SIMDU.scala 565:56 568:32]
  wire  _GEN_3180 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2452 : _GEN_1776; // @[SIMDU.scala 565:56]
  wire  _GEN_3181 = PMDU1_io_in_ready & ~match_operator_3 ? _GEN_2453 : _GEN_1777; // @[SIMDU.scala 565:56]
  wire  _GEN_3182 = PMDU0_io_in_ready & ~match_operator_2 | _GEN_1959; // @[SIMDU.scala 560:50 561:24]
  wire  _GEN_3361 = PMDU0_io_in_ready & ~match_operator_2 ? _GEN_2452 : _GEN_3180; // @[SIMDU.scala 560:50]
  wire  _GEN_3362 = PMDU0_io_in_ready & ~match_operator_2 ? _GEN_2453 : _GEN_3181; // @[SIMDU.scala 560:50]
  wire  _GEN_3363 = PMDU0_io_in_ready & ~match_operator_2 ? _GEN_2139 : _GEN_3001; // @[SIMDU.scala 560:50]
  wire  _GEN_3721 = _GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c) ? _GEN_3361 : _GEN_1776; // @[SIMDU.scala 559:142]
  wire  _GEN_3722 = _GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c) ? _GEN_3362 : _GEN_1777; // @[SIMDU.scala 559:142]
  wire  _T_66 = PALU0_io_out_bits_DecodeOut_InstNo <= PALU1_io_out_bits_DecodeOut_InstNo &
    PALU0_io_out_bits_DecodeOut_InstFlag == PALU1_io_out_bits_DecodeOut_InstFlag | PALU0_io_out_bits_DecodeOut_InstNo >
    PALU1_io_out_bits_DecodeOut_InstNo & PALU0_io_out_bits_DecodeOut_InstFlag != PALU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 450:101]
  wire  _T_67 = _T_66 ? 1'h0 : 1'h1; // @[SIMDU.scala 598:66]
  wire  winner0 = PALU0_io_out_valid ? PALU1_io_out_valid & _T_67 : 1'h1; // @[SIMDU.scala 598:20]
  wire  _T_75 = PMDU0_io_out_bits_DecodeOut_InstNo <= PMDU1_io_out_bits_DecodeOut_InstNo &
    PMDU0_io_out_bits_DecodeOut_InstFlag == PMDU1_io_out_bits_DecodeOut_InstFlag | PMDU0_io_out_bits_DecodeOut_InstNo >
    PMDU1_io_out_bits_DecodeOut_InstNo & PMDU0_io_out_bits_DecodeOut_InstFlag != PMDU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 450:101]
  wire [1:0] _T_76 = _T_75 ? 2'h2 : 2'h3; // @[SIMDU.scala 599:66]
  wire [1:0] _T_77 = PMDU1_io_out_valid ? _T_76 : 2'h2; // @[SIMDU.scala 599:43]
  wire [1:0] winner1 = PMDU0_io_out_valid ? _T_77 : 2'h3; // @[SIMDU.scala 599:20]
  wire  _T_78 = ~winner0; // @[SIMDU.scala 600:29]
  wire [4:0] InstNo0 = ~winner0 ? PALU0_io_out_bits_DecodeOut_InstNo : PALU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 600:20]
  wire  _T_79 = winner1 == 2'h2; // @[SIMDU.scala 601:29]
  wire [4:0] InstNo1 = winner1 == 2'h2 ? PMDU0_io_out_bits_DecodeOut_InstNo : PMDU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 601:20]
  wire  InstFlag0 = _T_78 ? PALU0_io_out_bits_DecodeOut_InstFlag : PALU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 602:22]
  wire  InstFlag1 = _T_79 ? PMDU0_io_out_bits_DecodeOut_InstFlag : PMDU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 603:22]
  wire  outvalid0 = _T_78 ? PALU0_io_out_valid : PALU1_io_out_valid; // @[SIMDU.scala 604:22]
  wire  outvalid1 = _T_79 ? PMDU0_io_out_valid : PMDU1_io_out_valid; // @[SIMDU.scala 605:22]
  wire  _T_90 = InstNo0 <= InstNo1 & InstFlag0 == InstFlag1 | InstNo0 > InstNo1 & InstFlag0 != InstFlag1; // @[SIMDU.scala 450:101]
  wire [1:0] _T_91 = _T_90 ? {{1'd0}, winner0} : winner1; // @[SIMDU.scala 606:46]
  wire [1:0] _T_92 = outvalid1 ? _T_91 : {{1'd0}, winner0}; // @[SIMDU.scala 606:32]
  wire [1:0] king = outvalid0 ? _T_92 : winner1; // @[SIMDU.scala 606:18]
  wire [1:0] _GEN_5054 = {{1'd0}, winner0}; // @[SIMDU.scala 607:24]
  wire  _T_93 = king == _GEN_5054; // @[SIMDU.scala 607:24]
  wire [1:0] queen0 = king == _GEN_5054 ? winner1 : {{1'd0}, winner0}; // @[SIMDU.scala 607:18]
  wire  _T_95 = king == 2'h0; // @[SIMDU.scala 608:45]
  wire  _T_97 = king == 2'h2; // @[SIMDU.scala 608:71]
  wire [1:0] _T_98 = king == 2'h2 ? 2'h3 : 2'h2; // @[SIMDU.scala 608:65]
  wire [1:0] queen1 = _T_93 ? {{1'd0}, king == 2'h0} : _T_98; // @[SIMDU.scala 608:18]
  wire  _T_99 = queen0 == 2'h0; // @[SIMDU.scala 609:28]
  wire  _T_100 = queen0 == 2'h1; // @[SIMDU.scala 609:82]
  wire  _T_101 = queen0 == 2'h2; // @[SIMDU.scala 609:136]
  wire [4:0] _T_102 = queen0 == 2'h2 ? PMDU0_io_out_bits_DecodeOut_InstNo : PMDU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 609:128]
  wire [4:0] _T_103 = queen0 == 2'h1 ? PALU1_io_out_bits_DecodeOut_InstNo : _T_102; // @[SIMDU.scala 609:74]
  wire [4:0] InstNo2 = queen0 == 2'h0 ? PALU0_io_out_bits_DecodeOut_InstNo : _T_103; // @[SIMDU.scala 609:20]
  wire  _T_104 = queen1 == 2'h0; // @[SIMDU.scala 610:28]
  wire  _T_105 = queen1 == 2'h1; // @[SIMDU.scala 610:82]
  wire  _T_106 = queen1 == 2'h2; // @[SIMDU.scala 610:136]
  wire [4:0] _T_107 = queen1 == 2'h2 ? PMDU0_io_out_bits_DecodeOut_InstNo : PMDU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 610:128]
  wire [4:0] _T_108 = queen1 == 2'h1 ? PALU1_io_out_bits_DecodeOut_InstNo : _T_107; // @[SIMDU.scala 610:74]
  wire [4:0] InstNo3 = queen1 == 2'h0 ? PALU0_io_out_bits_DecodeOut_InstNo : _T_108; // @[SIMDU.scala 610:20]
  wire  _T_112 = _T_101 ? PMDU0_io_out_bits_DecodeOut_InstFlag : PMDU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 611:134]
  wire  _T_113 = _T_100 ? PALU1_io_out_bits_DecodeOut_InstFlag : _T_112; // @[SIMDU.scala 611:78]
  wire  InstFlag2 = _T_99 ? PALU0_io_out_bits_DecodeOut_InstFlag : _T_113; // @[SIMDU.scala 611:22]
  wire  _T_117 = _T_106 ? PMDU0_io_out_bits_DecodeOut_InstFlag : PMDU1_io_out_bits_DecodeOut_InstFlag; // @[SIMDU.scala 612:134]
  wire  _T_118 = _T_105 ? PALU1_io_out_bits_DecodeOut_InstFlag : _T_117; // @[SIMDU.scala 612:78]
  wire  InstFlag3 = _T_104 ? PALU0_io_out_bits_DecodeOut_InstFlag : _T_118; // @[SIMDU.scala 612:22]
  wire  _T_122 = _T_101 ? PMDU0_io_out_valid : PMDU1_io_out_valid; // @[SIMDU.scala 613:98]
  wire  _T_123 = _T_100 ? PALU1_io_out_valid : _T_122; // @[SIMDU.scala 613:60]
  wire  outvalid2 = _T_99 ? PALU0_io_out_valid : _T_123; // @[SIMDU.scala 613:22]
  wire  _T_127 = _T_106 ? PMDU0_io_out_valid : PMDU1_io_out_valid; // @[SIMDU.scala 614:98]
  wire  _T_128 = _T_105 ? PALU1_io_out_valid : _T_127; // @[SIMDU.scala 614:60]
  wire  outvalid3 = _T_104 ? PALU0_io_out_valid : _T_128; // @[SIMDU.scala 614:22]
  wire  _T_135 = InstNo2 <= InstNo3 & InstFlag2 == InstFlag3 | InstNo2 > InstNo3 & InstFlag2 != InstFlag3; // @[SIMDU.scala 450:101]
  wire [1:0] _T_136 = _T_135 ? queen0 : queen1; // @[SIMDU.scala 615:46]
  wire [1:0] _T_137 = outvalid3 ? _T_136 : queen0; // @[SIMDU.scala 615:32]
  wire [1:0] queen = outvalid2 ? _T_137 : queen1; // @[SIMDU.scala 615:18]
  wire [63:0] _GEN_4624 = _T_97 ? PMDU0_io_out_bits_result : PMDU1_io_out_bits_result; // @[SIMDU.scala 627:27 628:20 633:20]
  wire [4:0] _GEN_4626 = _T_97 ? PMDU0_io_out_bits_DecodeOut_InstNo : PMDU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 627:27 629:20 634:20]
  wire  _GEN_4627 = _T_97 ? PMDU0_io_out_bits_DecodeOut_pext_OV : PMDU1_io_out_bits_DecodeOut_pext_OV; // @[SIMDU.scala 627:27 629:20 634:20]
  wire [4:0] _GEN_4639 = _T_97 ? PMDU0_io_out_bits_DecodeOut_ctrl_rfDest : PMDU1_io_out_bits_DecodeOut_ctrl_rfDest; // @[SIMDU.scala 627:27 629:20 634:20]
  wire  _GEN_4640 = _T_97 ? PMDU0_io_out_bits_DecodeOut_ctrl_rfWen : PMDU1_io_out_bits_DecodeOut_ctrl_rfWen; // @[SIMDU.scala 627:27 629:20 634:20]
  wire [63:0] _GEN_4653 = _T_97 ? PMDU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id :
    PMDU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id; // @[SIMDU.scala 627:27 629:20 634:20]
  wire [38:0] _GEN_4689 = _T_97 ? PMDU0_io_out_bits_DecodeOut_cf_pc : PMDU1_io_out_bits_DecodeOut_cf_pc; // @[SIMDU.scala 627:27 629:20 634:20]
  wire  _GEN_4691 = _T_97 ? PMDU0_io_out_valid : PMDU1_io_out_valid; // @[SIMDU.scala 627:27 630:20 635:20]
  wire  _GEN_4692 = _T_97 & io_out_0_ready; // @[SIMDU.scala 469:22 627:27 631:24]
  wire  _GEN_4693 = _T_97 ? 1'h0 : io_out_0_ready; // @[SIMDU.scala 471:22 627:27 636:24]
  wire [63:0] _GEN_4694 = king == 2'h1 ? PALU1_io_out_bits_result : _GEN_4624; // @[SIMDU.scala 622:27 623:20]
  wire [4:0] _GEN_4696 = king == 2'h1 ? PALU1_io_out_bits_DecodeOut_InstNo : _GEN_4626; // @[SIMDU.scala 622:27 624:20]
  wire  _GEN_4697 = king == 2'h1 ? PALU1_io_out_bits_DecodeOut_pext_OV : _GEN_4627; // @[SIMDU.scala 622:27 624:20]
  wire [4:0] _GEN_4709 = king == 2'h1 ? PALU1_io_out_bits_DecodeOut_ctrl_rfDest : _GEN_4639; // @[SIMDU.scala 622:27 624:20]
  wire  _GEN_4710 = king == 2'h1 ? PALU1_io_out_bits_DecodeOut_ctrl_rfWen : _GEN_4640; // @[SIMDU.scala 622:27 624:20]
  wire [63:0] _GEN_4723 = king == 2'h1 ? PALU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id : _GEN_4653; // @[SIMDU.scala 622:27 624:20]
  wire [38:0] _GEN_4759 = king == 2'h1 ? PALU1_io_out_bits_DecodeOut_cf_pc : _GEN_4689; // @[SIMDU.scala 622:27 624:20]
  wire  _GEN_4761 = king == 2'h1 ? PALU1_io_out_valid : _GEN_4691; // @[SIMDU.scala 622:27 625:20]
  wire  _GEN_4762 = king == 2'h1 & io_out_0_ready; // @[SIMDU.scala 470:22 622:27 626:24]
  wire  _GEN_4763 = king == 2'h1 ? 1'h0 : _GEN_4692; // @[SIMDU.scala 469:22 622:27]
  wire  _GEN_4764 = king == 2'h1 ? 1'h0 : _GEN_4693; // @[SIMDU.scala 471:22 622:27]
  wire  _GEN_4833 = _T_95 & io_out_0_ready; // @[SIMDU.scala 617:21 468:22 621:24]
  wire  _GEN_4834 = _T_95 ? 1'h0 : _GEN_4762; // @[SIMDU.scala 617:21 470:22]
  wire  _GEN_4835 = _T_95 ? 1'h0 : _GEN_4763; // @[SIMDU.scala 617:21 469:22]
  wire  _GEN_4836 = _T_95 ? 1'h0 : _GEN_4764; // @[SIMDU.scala 617:21 471:22]
  wire [63:0] _GEN_4837 = queen == 2'h2 ? PMDU0_io_out_bits_result : PMDU1_io_out_bits_result; // @[SIMDU.scala 648:28 649:20 654:20]
  wire [4:0] _GEN_4839 = queen == 2'h2 ? PMDU0_io_out_bits_DecodeOut_InstNo : PMDU1_io_out_bits_DecodeOut_InstNo; // @[SIMDU.scala 648:28 650:20 655:20]
  wire  _GEN_4840 = queen == 2'h2 ? PMDU0_io_out_bits_DecodeOut_pext_OV : PMDU1_io_out_bits_DecodeOut_pext_OV; // @[SIMDU.scala 648:28 650:20 655:20]
  wire [4:0] _GEN_4852 = queen == 2'h2 ? PMDU0_io_out_bits_DecodeOut_ctrl_rfDest :
    PMDU1_io_out_bits_DecodeOut_ctrl_rfDest; // @[SIMDU.scala 648:28 650:20 655:20]
  wire  _GEN_4853 = queen == 2'h2 ? PMDU0_io_out_bits_DecodeOut_ctrl_rfWen : PMDU1_io_out_bits_DecodeOut_ctrl_rfWen; // @[SIMDU.scala 648:28 650:20 655:20]
  wire [63:0] _GEN_4866 = queen == 2'h2 ? PMDU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id :
    PMDU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id; // @[SIMDU.scala 648:28 650:20 655:20]
  wire [38:0] _GEN_4902 = queen == 2'h2 ? PMDU0_io_out_bits_DecodeOut_cf_pc : PMDU1_io_out_bits_DecodeOut_cf_pc; // @[SIMDU.scala 648:28 650:20 655:20]
  wire  _GEN_4904 = queen == 2'h2 ? PMDU0_io_out_valid : PMDU1_io_out_valid; // @[SIMDU.scala 648:28 651:20 656:20]
  wire  _GEN_4905 = queen == 2'h2 ? io_out_1_ready : _GEN_4835; // @[SIMDU.scala 648:28 652:24]
  wire  _GEN_4906 = queen == 2'h2 ? _GEN_4836 : io_out_1_ready; // @[SIMDU.scala 648:28 657:24]
  wire [63:0] _GEN_4907 = queen == 2'h1 ? PALU1_io_out_bits_result : _GEN_4837; // @[SIMDU.scala 643:28 644:20]
  wire [4:0] _GEN_4909 = queen == 2'h1 ? PALU1_io_out_bits_DecodeOut_InstNo : _GEN_4839; // @[SIMDU.scala 643:28 645:20]
  wire  _GEN_4910 = queen == 2'h1 ? PALU1_io_out_bits_DecodeOut_pext_OV : _GEN_4840; // @[SIMDU.scala 643:28 645:20]
  wire [4:0] _GEN_4922 = queen == 2'h1 ? PALU1_io_out_bits_DecodeOut_ctrl_rfDest : _GEN_4852; // @[SIMDU.scala 643:28 645:20]
  wire  _GEN_4923 = queen == 2'h1 ? PALU1_io_out_bits_DecodeOut_ctrl_rfWen : _GEN_4853; // @[SIMDU.scala 643:28 645:20]
  wire [63:0] _GEN_4936 = queen == 2'h1 ? PALU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id : _GEN_4866; // @[SIMDU.scala 643:28 645:20]
  wire [38:0] _GEN_4972 = queen == 2'h1 ? PALU1_io_out_bits_DecodeOut_cf_pc : _GEN_4902; // @[SIMDU.scala 643:28 645:20]
  wire  _GEN_4974 = queen == 2'h1 ? PALU1_io_out_valid : _GEN_4904; // @[SIMDU.scala 643:28 646:20]
  wire  _GEN_4975 = queen == 2'h1 ? io_out_1_ready : _GEN_4834; // @[SIMDU.scala 643:28 647:24]
  wire  _GEN_4976 = queen == 2'h1 ? _GEN_4835 : _GEN_4905; // @[SIMDU.scala 643:28]
  wire  _GEN_4977 = queen == 2'h1 ? _GEN_4836 : _GEN_4906; // @[SIMDU.scala 643:28]
  PALU PALU0 ( // @[SIMDU.scala 451:21]
    .io_in_ready(PALU0_io_in_ready),
    .io_in_valid(PALU0_io_in_valid),
    .io_in_bits_DecodeIn_cf_pc(PALU0_io_in_bits_DecodeIn_cf_pc),
    .io_in_bits_DecodeIn_cf_runahead_checkpoint_id(PALU0_io_in_bits_DecodeIn_cf_runahead_checkpoint_id),
    .io_in_bits_DecodeIn_ctrl_fuOpType(PALU0_io_in_bits_DecodeIn_ctrl_fuOpType),
    .io_in_bits_DecodeIn_ctrl_funct3(PALU0_io_in_bits_DecodeIn_ctrl_funct3),
    .io_in_bits_DecodeIn_ctrl_func24(PALU0_io_in_bits_DecodeIn_ctrl_func24),
    .io_in_bits_DecodeIn_ctrl_rfWen(PALU0_io_in_bits_DecodeIn_ctrl_rfWen),
    .io_in_bits_DecodeIn_ctrl_rfDest(PALU0_io_in_bits_DecodeIn_ctrl_rfDest),
    .io_in_bits_DecodeIn_data_src1(PALU0_io_in_bits_DecodeIn_data_src1),
    .io_in_bits_DecodeIn_data_src2(PALU0_io_in_bits_DecodeIn_data_src2),
    .io_in_bits_DecodeIn_data_src3(PALU0_io_in_bits_DecodeIn_data_src3),
    .io_in_bits_DecodeIn_InstNo(PALU0_io_in_bits_DecodeIn_InstNo),
    .io_in_bits_DecodeIn_InstFlag(PALU0_io_in_bits_DecodeIn_InstFlag),
    .io_in_bits_Pctrl_isAdd_64(PALU0_io_in_bits_Pctrl_isAdd_64),
    .io_in_bits_Pctrl_isAdd_32(PALU0_io_in_bits_Pctrl_isAdd_32),
    .io_in_bits_Pctrl_isAdd_16(PALU0_io_in_bits_Pctrl_isAdd_16),
    .io_in_bits_Pctrl_isAdd_8(PALU0_io_in_bits_Pctrl_isAdd_8),
    .io_in_bits_Pctrl_isAdd_Q15(PALU0_io_in_bits_Pctrl_isAdd_Q15),
    .io_in_bits_Pctrl_isAdd_Q31(PALU0_io_in_bits_Pctrl_isAdd_Q31),
    .io_in_bits_Pctrl_isAdd_C31(PALU0_io_in_bits_Pctrl_isAdd_C31),
    .io_in_bits_Pctrl_isAve(PALU0_io_in_bits_Pctrl_isAve),
    .io_in_bits_Pctrl_isSub_64(PALU0_io_in_bits_Pctrl_isSub_64),
    .io_in_bits_Pctrl_isSub_32(PALU0_io_in_bits_Pctrl_isSub_32),
    .io_in_bits_Pctrl_isSub_16(PALU0_io_in_bits_Pctrl_isSub_16),
    .io_in_bits_Pctrl_isSub_8(PALU0_io_in_bits_Pctrl_isSub_8),
    .io_in_bits_Pctrl_isSub_Q15(PALU0_io_in_bits_Pctrl_isSub_Q15),
    .io_in_bits_Pctrl_isSub_Q31(PALU0_io_in_bits_Pctrl_isSub_Q31),
    .io_in_bits_Pctrl_isSub_C31(PALU0_io_in_bits_Pctrl_isSub_C31),
    .io_in_bits_Pctrl_isCras_16(PALU0_io_in_bits_Pctrl_isCras_16),
    .io_in_bits_Pctrl_isCrsa_16(PALU0_io_in_bits_Pctrl_isCrsa_16),
    .io_in_bits_Pctrl_isCras_32(PALU0_io_in_bits_Pctrl_isCras_32),
    .io_in_bits_Pctrl_isCrsa_32(PALU0_io_in_bits_Pctrl_isCrsa_32),
    .io_in_bits_Pctrl_isStas_16(PALU0_io_in_bits_Pctrl_isStas_16),
    .io_in_bits_Pctrl_isStsa_16(PALU0_io_in_bits_Pctrl_isStsa_16),
    .io_in_bits_Pctrl_isStas_32(PALU0_io_in_bits_Pctrl_isStas_32),
    .io_in_bits_Pctrl_isStsa_32(PALU0_io_in_bits_Pctrl_isStsa_32),
    .io_in_bits_Pctrl_isComp_16(PALU0_io_in_bits_Pctrl_isComp_16),
    .io_in_bits_Pctrl_isComp_8(PALU0_io_in_bits_Pctrl_isComp_8),
    .io_in_bits_Pctrl_isCompare(PALU0_io_in_bits_Pctrl_isCompare),
    .io_in_bits_Pctrl_isMaxMin_16(PALU0_io_in_bits_Pctrl_isMaxMin_16),
    .io_in_bits_Pctrl_isMaxMin_8(PALU0_io_in_bits_Pctrl_isMaxMin_8),
    .io_in_bits_Pctrl_isMaxMin_XLEN(PALU0_io_in_bits_Pctrl_isMaxMin_XLEN),
    .io_in_bits_Pctrl_isMaxMin_32(PALU0_io_in_bits_Pctrl_isMaxMin_32),
    .io_in_bits_Pctrl_isMaxMin(PALU0_io_in_bits_Pctrl_isMaxMin),
    .io_in_bits_Pctrl_isPbs(PALU0_io_in_bits_Pctrl_isPbs),
    .io_in_bits_Pctrl_isRs_16(PALU0_io_in_bits_Pctrl_isRs_16),
    .io_in_bits_Pctrl_isLs_16(PALU0_io_in_bits_Pctrl_isLs_16),
    .io_in_bits_Pctrl_isLR_16(PALU0_io_in_bits_Pctrl_isLR_16),
    .io_in_bits_Pctrl_isRs_8(PALU0_io_in_bits_Pctrl_isRs_8),
    .io_in_bits_Pctrl_isLs_8(PALU0_io_in_bits_Pctrl_isLs_8),
    .io_in_bits_Pctrl_isLR_8(PALU0_io_in_bits_Pctrl_isLR_8),
    .io_in_bits_Pctrl_isRs_32(PALU0_io_in_bits_Pctrl_isRs_32),
    .io_in_bits_Pctrl_isLs_32(PALU0_io_in_bits_Pctrl_isLs_32),
    .io_in_bits_Pctrl_isLR_32(PALU0_io_in_bits_Pctrl_isLR_32),
    .io_in_bits_Pctrl_isLR_Q31(PALU0_io_in_bits_Pctrl_isLR_Q31),
    .io_in_bits_Pctrl_isLs_Q31(PALU0_io_in_bits_Pctrl_isLs_Q31),
    .io_in_bits_Pctrl_isRs_XLEN(PALU0_io_in_bits_Pctrl_isRs_XLEN),
    .io_in_bits_Pctrl_isSRAIWU(PALU0_io_in_bits_Pctrl_isSRAIWU),
    .io_in_bits_Pctrl_isFSRW(PALU0_io_in_bits_Pctrl_isFSRW),
    .io_in_bits_Pctrl_isWext(PALU0_io_in_bits_Pctrl_isWext),
    .io_in_bits_Pctrl_isShifter(PALU0_io_in_bits_Pctrl_isShifter),
    .io_in_bits_Pctrl_isClip_16(PALU0_io_in_bits_Pctrl_isClip_16),
    .io_in_bits_Pctrl_isClip_8(PALU0_io_in_bits_Pctrl_isClip_8),
    .io_in_bits_Pctrl_isclip_32(PALU0_io_in_bits_Pctrl_isclip_32),
    .io_in_bits_Pctrl_isClip(PALU0_io_in_bits_Pctrl_isClip),
    .io_in_bits_Pctrl_isSat_16(PALU0_io_in_bits_Pctrl_isSat_16),
    .io_in_bits_Pctrl_isSat_8(PALU0_io_in_bits_Pctrl_isSat_8),
    .io_in_bits_Pctrl_isSat_32(PALU0_io_in_bits_Pctrl_isSat_32),
    .io_in_bits_Pctrl_isSat_W(PALU0_io_in_bits_Pctrl_isSat_W),
    .io_in_bits_Pctrl_isSat(PALU0_io_in_bits_Pctrl_isSat),
    .io_in_bits_Pctrl_isCnt_16(PALU0_io_in_bits_Pctrl_isCnt_16),
    .io_in_bits_Pctrl_isCnt_8(PALU0_io_in_bits_Pctrl_isCnt_8),
    .io_in_bits_Pctrl_isCnt_32(PALU0_io_in_bits_Pctrl_isCnt_32),
    .io_in_bits_Pctrl_isCnt(PALU0_io_in_bits_Pctrl_isCnt),
    .io_in_bits_Pctrl_isSwap_16(PALU0_io_in_bits_Pctrl_isSwap_16),
    .io_in_bits_Pctrl_isSwap_8(PALU0_io_in_bits_Pctrl_isSwap_8),
    .io_in_bits_Pctrl_isSwap(PALU0_io_in_bits_Pctrl_isSwap),
    .io_in_bits_Pctrl_isUnpack(PALU0_io_in_bits_Pctrl_isUnpack),
    .io_in_bits_Pctrl_isBitrev(PALU0_io_in_bits_Pctrl_isBitrev),
    .io_in_bits_Pctrl_isCmix(PALU0_io_in_bits_Pctrl_isCmix),
    .io_in_bits_Pctrl_isInsertb(PALU0_io_in_bits_Pctrl_isInsertb),
    .io_in_bits_Pctrl_isPackbb(PALU0_io_in_bits_Pctrl_isPackbb),
    .io_in_bits_Pctrl_isPackbt(PALU0_io_in_bits_Pctrl_isPackbt),
    .io_in_bits_Pctrl_isPacktb(PALU0_io_in_bits_Pctrl_isPacktb),
    .io_in_bits_Pctrl_isPacktt(PALU0_io_in_bits_Pctrl_isPacktt),
    .io_in_bits_Pctrl_isPack(PALU0_io_in_bits_Pctrl_isPack),
    .io_in_bits_Pctrl_isSub(PALU0_io_in_bits_Pctrl_isSub),
    .io_in_bits_Pctrl_isAdder(PALU0_io_in_bits_Pctrl_isAdder),
    .io_in_bits_Pctrl_SrcSigned(PALU0_io_in_bits_Pctrl_SrcSigned),
    .io_in_bits_Pctrl_Saturating(PALU0_io_in_bits_Pctrl_Saturating),
    .io_in_bits_Pctrl_Translation(PALU0_io_in_bits_Pctrl_Translation),
    .io_in_bits_Pctrl_LessEqual(PALU0_io_in_bits_Pctrl_LessEqual),
    .io_in_bits_Pctrl_LessThan(PALU0_io_in_bits_Pctrl_LessThan),
    .io_in_bits_Pctrl_adderRes_ori(PALU0_io_in_bits_Pctrl_adderRes_ori),
    .io_in_bits_Pctrl_adderRes(PALU0_io_in_bits_Pctrl_adderRes),
    .io_in_bits_Pctrl_adderRes_ori_drophighestbit(PALU0_io_in_bits_Pctrl_adderRes_ori_drophighestbit),
    .io_in_bits_Pctrl_Round(PALU0_io_in_bits_Pctrl_Round),
    .io_in_bits_Pctrl_ShiftSigned(PALU0_io_in_bits_Pctrl_ShiftSigned),
    .io_in_bits_Pctrl_Arithmetic(PALU0_io_in_bits_Pctrl_Arithmetic),
    .io_out_ready(PALU0_io_out_ready),
    .io_out_valid(PALU0_io_out_valid),
    .io_out_bits_result(PALU0_io_out_bits_result),
    .io_out_bits_DecodeOut_cf_pc(PALU0_io_out_bits_DecodeOut_cf_pc),
    .io_out_bits_DecodeOut_cf_runahead_checkpoint_id(PALU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id),
    .io_out_bits_DecodeOut_ctrl_rfWen(PALU0_io_out_bits_DecodeOut_ctrl_rfWen),
    .io_out_bits_DecodeOut_ctrl_rfDest(PALU0_io_out_bits_DecodeOut_ctrl_rfDest),
    .io_out_bits_DecodeOut_pext_OV(PALU0_io_out_bits_DecodeOut_pext_OV),
    .io_out_bits_DecodeOut_InstNo(PALU0_io_out_bits_DecodeOut_InstNo),
    .io_out_bits_DecodeOut_InstFlag(PALU0_io_out_bits_DecodeOut_InstFlag)
  );
  PMDU PMDU0 ( // @[SIMDU.scala 452:21]
    .io_in_ready(PMDU0_io_in_ready),
    .io_in_valid(PMDU0_io_in_valid),
    .io_in_bits_DecodeIn_cf_pc(PMDU0_io_in_bits_DecodeIn_cf_pc),
    .io_in_bits_DecodeIn_cf_runahead_checkpoint_id(PMDU0_io_in_bits_DecodeIn_cf_runahead_checkpoint_id),
    .io_in_bits_DecodeIn_ctrl_fuOpType(PMDU0_io_in_bits_DecodeIn_ctrl_fuOpType),
    .io_in_bits_DecodeIn_ctrl_rfWen(PMDU0_io_in_bits_DecodeIn_ctrl_rfWen),
    .io_in_bits_DecodeIn_ctrl_rfDest(PMDU0_io_in_bits_DecodeIn_ctrl_rfDest),
    .io_in_bits_DecodeIn_data_src1(PMDU0_io_in_bits_DecodeIn_data_src1),
    .io_in_bits_DecodeIn_data_src2(PMDU0_io_in_bits_DecodeIn_data_src2),
    .io_in_bits_DecodeIn_data_src3(PMDU0_io_in_bits_DecodeIn_data_src3),
    .io_in_bits_DecodeIn_InstNo(PMDU0_io_in_bits_DecodeIn_InstNo),
    .io_in_bits_DecodeIn_InstFlag(PMDU0_io_in_bits_DecodeIn_InstFlag),
    .io_in_bits_Pctrl_isMul_16(PMDU0_io_in_bits_Pctrl_isMul_16),
    .io_in_bits_Pctrl_isMul_8(PMDU0_io_in_bits_Pctrl_isMul_8),
    .io_in_bits_Pctrl_isMSW_3232(PMDU0_io_in_bits_Pctrl_isMSW_3232),
    .io_in_bits_Pctrl_isMSW_3216(PMDU0_io_in_bits_Pctrl_isMSW_3216),
    .io_in_bits_Pctrl_isS1632(PMDU0_io_in_bits_Pctrl_isS1632),
    .io_in_bits_Pctrl_isS1664(PMDU0_io_in_bits_Pctrl_isS1664),
    .io_in_bits_Pctrl_is832(PMDU0_io_in_bits_Pctrl_is832),
    .io_in_bits_Pctrl_is3264(PMDU0_io_in_bits_Pctrl_is3264),
    .io_in_bits_Pctrl_is1664(PMDU0_io_in_bits_Pctrl_is1664),
    .io_in_bits_Pctrl_isQ15orQ31(PMDU0_io_in_bits_Pctrl_isQ15orQ31),
    .io_in_bits_Pctrl_isC31(PMDU0_io_in_bits_Pctrl_isC31),
    .io_in_bits_Pctrl_isQ15_64ONLY(PMDU0_io_in_bits_Pctrl_isQ15_64ONLY),
    .io_in_bits_Pctrl_isQ63_64ONLY(PMDU0_io_in_bits_Pctrl_isQ63_64ONLY),
    .io_in_bits_Pctrl_isMul_32_64ONLY(PMDU0_io_in_bits_Pctrl_isMul_32_64ONLY),
    .io_in_bits_Pctrl_isPMA_64ONLY(PMDU0_io_in_bits_Pctrl_isPMA_64ONLY),
    .io_in_bits_Pctrl_mulres9_0(PMDU0_io_in_bits_Pctrl_mulres9_0),
    .io_in_bits_Pctrl_mulres9_1(PMDU0_io_in_bits_Pctrl_mulres9_1),
    .io_in_bits_Pctrl_mulres9_2(PMDU0_io_in_bits_Pctrl_mulres9_2),
    .io_in_bits_Pctrl_mulres9_3(PMDU0_io_in_bits_Pctrl_mulres9_3),
    .io_in_bits_Pctrl_mulres17_0(PMDU0_io_in_bits_Pctrl_mulres17_0),
    .io_in_bits_Pctrl_mulres17_1(PMDU0_io_in_bits_Pctrl_mulres17_1),
    .io_in_bits_Pctrl_mulres33_0(PMDU0_io_in_bits_Pctrl_mulres33_0),
    .io_in_bits_Pctrl_mulres65_0(PMDU0_io_in_bits_Pctrl_mulres65_0),
    .io_out_ready(PMDU0_io_out_ready),
    .io_out_valid(PMDU0_io_out_valid),
    .io_out_bits_result(PMDU0_io_out_bits_result),
    .io_out_bits_DecodeOut_cf_pc(PMDU0_io_out_bits_DecodeOut_cf_pc),
    .io_out_bits_DecodeOut_cf_runahead_checkpoint_id(PMDU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id),
    .io_out_bits_DecodeOut_ctrl_fuOpType(PMDU0_io_out_bits_DecodeOut_ctrl_fuOpType),
    .io_out_bits_DecodeOut_ctrl_rfWen(PMDU0_io_out_bits_DecodeOut_ctrl_rfWen),
    .io_out_bits_DecodeOut_ctrl_rfDest(PMDU0_io_out_bits_DecodeOut_ctrl_rfDest),
    .io_out_bits_DecodeOut_data_src1(PMDU0_io_out_bits_DecodeOut_data_src1),
    .io_out_bits_DecodeOut_data_src2(PMDU0_io_out_bits_DecodeOut_data_src2),
    .io_out_bits_DecodeOut_data_src3(PMDU0_io_out_bits_DecodeOut_data_src3),
    .io_out_bits_DecodeOut_pext_OV(PMDU0_io_out_bits_DecodeOut_pext_OV),
    .io_out_bits_DecodeOut_InstNo(PMDU0_io_out_bits_DecodeOut_InstNo),
    .io_out_bits_DecodeOut_InstFlag(PMDU0_io_out_bits_DecodeOut_InstFlag),
    .io_FirstStageFire(PMDU0_io_FirstStageFire)
  );
  PALU_1 PALU1 ( // @[SIMDU.scala 453:21]
    .io_in_ready(PALU1_io_in_ready),
    .io_in_valid(PALU1_io_in_valid),
    .io_in_bits_DecodeIn_cf_pc(PALU1_io_in_bits_DecodeIn_cf_pc),
    .io_in_bits_DecodeIn_cf_runahead_checkpoint_id(PALU1_io_in_bits_DecodeIn_cf_runahead_checkpoint_id),
    .io_in_bits_DecodeIn_ctrl_fuOpType(PALU1_io_in_bits_DecodeIn_ctrl_fuOpType),
    .io_in_bits_DecodeIn_ctrl_funct3(PALU1_io_in_bits_DecodeIn_ctrl_funct3),
    .io_in_bits_DecodeIn_ctrl_func24(PALU1_io_in_bits_DecodeIn_ctrl_func24),
    .io_in_bits_DecodeIn_ctrl_rfWen(PALU1_io_in_bits_DecodeIn_ctrl_rfWen),
    .io_in_bits_DecodeIn_ctrl_rfDest(PALU1_io_in_bits_DecodeIn_ctrl_rfDest),
    .io_in_bits_DecodeIn_data_src1(PALU1_io_in_bits_DecodeIn_data_src1),
    .io_in_bits_DecodeIn_data_src2(PALU1_io_in_bits_DecodeIn_data_src2),
    .io_in_bits_DecodeIn_data_src3(PALU1_io_in_bits_DecodeIn_data_src3),
    .io_in_bits_DecodeIn_InstNo(PALU1_io_in_bits_DecodeIn_InstNo),
    .io_in_bits_DecodeIn_InstFlag(PALU1_io_in_bits_DecodeIn_InstFlag),
    .io_in_bits_Pctrl_isAdd_64(PALU1_io_in_bits_Pctrl_isAdd_64),
    .io_in_bits_Pctrl_isAdd_32(PALU1_io_in_bits_Pctrl_isAdd_32),
    .io_in_bits_Pctrl_isAdd_16(PALU1_io_in_bits_Pctrl_isAdd_16),
    .io_in_bits_Pctrl_isAdd_8(PALU1_io_in_bits_Pctrl_isAdd_8),
    .io_in_bits_Pctrl_isAdd_Q15(PALU1_io_in_bits_Pctrl_isAdd_Q15),
    .io_in_bits_Pctrl_isAdd_Q31(PALU1_io_in_bits_Pctrl_isAdd_Q31),
    .io_in_bits_Pctrl_isAdd_C31(PALU1_io_in_bits_Pctrl_isAdd_C31),
    .io_in_bits_Pctrl_isAve(PALU1_io_in_bits_Pctrl_isAve),
    .io_in_bits_Pctrl_isSub_64(PALU1_io_in_bits_Pctrl_isSub_64),
    .io_in_bits_Pctrl_isSub_32(PALU1_io_in_bits_Pctrl_isSub_32),
    .io_in_bits_Pctrl_isSub_16(PALU1_io_in_bits_Pctrl_isSub_16),
    .io_in_bits_Pctrl_isSub_8(PALU1_io_in_bits_Pctrl_isSub_8),
    .io_in_bits_Pctrl_isSub_Q15(PALU1_io_in_bits_Pctrl_isSub_Q15),
    .io_in_bits_Pctrl_isSub_Q31(PALU1_io_in_bits_Pctrl_isSub_Q31),
    .io_in_bits_Pctrl_isSub_C31(PALU1_io_in_bits_Pctrl_isSub_C31),
    .io_in_bits_Pctrl_isCras_16(PALU1_io_in_bits_Pctrl_isCras_16),
    .io_in_bits_Pctrl_isCrsa_16(PALU1_io_in_bits_Pctrl_isCrsa_16),
    .io_in_bits_Pctrl_isCras_32(PALU1_io_in_bits_Pctrl_isCras_32),
    .io_in_bits_Pctrl_isCrsa_32(PALU1_io_in_bits_Pctrl_isCrsa_32),
    .io_in_bits_Pctrl_isStas_16(PALU1_io_in_bits_Pctrl_isStas_16),
    .io_in_bits_Pctrl_isStsa_16(PALU1_io_in_bits_Pctrl_isStsa_16),
    .io_in_bits_Pctrl_isStas_32(PALU1_io_in_bits_Pctrl_isStas_32),
    .io_in_bits_Pctrl_isStsa_32(PALU1_io_in_bits_Pctrl_isStsa_32),
    .io_in_bits_Pctrl_isComp_16(PALU1_io_in_bits_Pctrl_isComp_16),
    .io_in_bits_Pctrl_isComp_8(PALU1_io_in_bits_Pctrl_isComp_8),
    .io_in_bits_Pctrl_isCompare(PALU1_io_in_bits_Pctrl_isCompare),
    .io_in_bits_Pctrl_isMaxMin_16(PALU1_io_in_bits_Pctrl_isMaxMin_16),
    .io_in_bits_Pctrl_isMaxMin_8(PALU1_io_in_bits_Pctrl_isMaxMin_8),
    .io_in_bits_Pctrl_isMaxMin_XLEN(PALU1_io_in_bits_Pctrl_isMaxMin_XLEN),
    .io_in_bits_Pctrl_isMaxMin_32(PALU1_io_in_bits_Pctrl_isMaxMin_32),
    .io_in_bits_Pctrl_isMaxMin(PALU1_io_in_bits_Pctrl_isMaxMin),
    .io_in_bits_Pctrl_isPbs(PALU1_io_in_bits_Pctrl_isPbs),
    .io_in_bits_Pctrl_isRs_16(PALU1_io_in_bits_Pctrl_isRs_16),
    .io_in_bits_Pctrl_isLs_16(PALU1_io_in_bits_Pctrl_isLs_16),
    .io_in_bits_Pctrl_isLR_16(PALU1_io_in_bits_Pctrl_isLR_16),
    .io_in_bits_Pctrl_isRs_8(PALU1_io_in_bits_Pctrl_isRs_8),
    .io_in_bits_Pctrl_isLs_8(PALU1_io_in_bits_Pctrl_isLs_8),
    .io_in_bits_Pctrl_isLR_8(PALU1_io_in_bits_Pctrl_isLR_8),
    .io_in_bits_Pctrl_isRs_32(PALU1_io_in_bits_Pctrl_isRs_32),
    .io_in_bits_Pctrl_isLs_32(PALU1_io_in_bits_Pctrl_isLs_32),
    .io_in_bits_Pctrl_isLR_32(PALU1_io_in_bits_Pctrl_isLR_32),
    .io_in_bits_Pctrl_isLR_Q31(PALU1_io_in_bits_Pctrl_isLR_Q31),
    .io_in_bits_Pctrl_isLs_Q31(PALU1_io_in_bits_Pctrl_isLs_Q31),
    .io_in_bits_Pctrl_isRs_XLEN(PALU1_io_in_bits_Pctrl_isRs_XLEN),
    .io_in_bits_Pctrl_isSRAIWU(PALU1_io_in_bits_Pctrl_isSRAIWU),
    .io_in_bits_Pctrl_isFSRW(PALU1_io_in_bits_Pctrl_isFSRW),
    .io_in_bits_Pctrl_isWext(PALU1_io_in_bits_Pctrl_isWext),
    .io_in_bits_Pctrl_isShifter(PALU1_io_in_bits_Pctrl_isShifter),
    .io_in_bits_Pctrl_isClip_16(PALU1_io_in_bits_Pctrl_isClip_16),
    .io_in_bits_Pctrl_isClip_8(PALU1_io_in_bits_Pctrl_isClip_8),
    .io_in_bits_Pctrl_isclip_32(PALU1_io_in_bits_Pctrl_isclip_32),
    .io_in_bits_Pctrl_isClip(PALU1_io_in_bits_Pctrl_isClip),
    .io_in_bits_Pctrl_isSat_16(PALU1_io_in_bits_Pctrl_isSat_16),
    .io_in_bits_Pctrl_isSat_8(PALU1_io_in_bits_Pctrl_isSat_8),
    .io_in_bits_Pctrl_isSat_32(PALU1_io_in_bits_Pctrl_isSat_32),
    .io_in_bits_Pctrl_isSat_W(PALU1_io_in_bits_Pctrl_isSat_W),
    .io_in_bits_Pctrl_isSat(PALU1_io_in_bits_Pctrl_isSat),
    .io_in_bits_Pctrl_isCnt_16(PALU1_io_in_bits_Pctrl_isCnt_16),
    .io_in_bits_Pctrl_isCnt_8(PALU1_io_in_bits_Pctrl_isCnt_8),
    .io_in_bits_Pctrl_isCnt_32(PALU1_io_in_bits_Pctrl_isCnt_32),
    .io_in_bits_Pctrl_isCnt(PALU1_io_in_bits_Pctrl_isCnt),
    .io_in_bits_Pctrl_isSwap_16(PALU1_io_in_bits_Pctrl_isSwap_16),
    .io_in_bits_Pctrl_isSwap_8(PALU1_io_in_bits_Pctrl_isSwap_8),
    .io_in_bits_Pctrl_isSwap(PALU1_io_in_bits_Pctrl_isSwap),
    .io_in_bits_Pctrl_isUnpack(PALU1_io_in_bits_Pctrl_isUnpack),
    .io_in_bits_Pctrl_isBitrev(PALU1_io_in_bits_Pctrl_isBitrev),
    .io_in_bits_Pctrl_isCmix(PALU1_io_in_bits_Pctrl_isCmix),
    .io_in_bits_Pctrl_isInsertb(PALU1_io_in_bits_Pctrl_isInsertb),
    .io_in_bits_Pctrl_isPackbb(PALU1_io_in_bits_Pctrl_isPackbb),
    .io_in_bits_Pctrl_isPackbt(PALU1_io_in_bits_Pctrl_isPackbt),
    .io_in_bits_Pctrl_isPacktb(PALU1_io_in_bits_Pctrl_isPacktb),
    .io_in_bits_Pctrl_isPacktt(PALU1_io_in_bits_Pctrl_isPacktt),
    .io_in_bits_Pctrl_isPack(PALU1_io_in_bits_Pctrl_isPack),
    .io_in_bits_Pctrl_isSub(PALU1_io_in_bits_Pctrl_isSub),
    .io_in_bits_Pctrl_isAdder(PALU1_io_in_bits_Pctrl_isAdder),
    .io_in_bits_Pctrl_SrcSigned(PALU1_io_in_bits_Pctrl_SrcSigned),
    .io_in_bits_Pctrl_Saturating(PALU1_io_in_bits_Pctrl_Saturating),
    .io_in_bits_Pctrl_Translation(PALU1_io_in_bits_Pctrl_Translation),
    .io_in_bits_Pctrl_LessEqual(PALU1_io_in_bits_Pctrl_LessEqual),
    .io_in_bits_Pctrl_LessThan(PALU1_io_in_bits_Pctrl_LessThan),
    .io_in_bits_Pctrl_adderRes_ori(PALU1_io_in_bits_Pctrl_adderRes_ori),
    .io_in_bits_Pctrl_adderRes(PALU1_io_in_bits_Pctrl_adderRes),
    .io_in_bits_Pctrl_adderRes_ori_drophighestbit(PALU1_io_in_bits_Pctrl_adderRes_ori_drophighestbit),
    .io_in_bits_Pctrl_Round(PALU1_io_in_bits_Pctrl_Round),
    .io_in_bits_Pctrl_ShiftSigned(PALU1_io_in_bits_Pctrl_ShiftSigned),
    .io_in_bits_Pctrl_Arithmetic(PALU1_io_in_bits_Pctrl_Arithmetic),
    .io_out_ready(PALU1_io_out_ready),
    .io_out_valid(PALU1_io_out_valid),
    .io_out_bits_result(PALU1_io_out_bits_result),
    .io_out_bits_DecodeOut_cf_pc(PALU1_io_out_bits_DecodeOut_cf_pc),
    .io_out_bits_DecodeOut_cf_runahead_checkpoint_id(PALU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id),
    .io_out_bits_DecodeOut_ctrl_rfWen(PALU1_io_out_bits_DecodeOut_ctrl_rfWen),
    .io_out_bits_DecodeOut_ctrl_rfDest(PALU1_io_out_bits_DecodeOut_ctrl_rfDest),
    .io_out_bits_DecodeOut_pext_OV(PALU1_io_out_bits_DecodeOut_pext_OV),
    .io_out_bits_DecodeOut_InstNo(PALU1_io_out_bits_DecodeOut_InstNo),
    .io_out_bits_DecodeOut_InstFlag(PALU1_io_out_bits_DecodeOut_InstFlag)
  );
  PMDU_1 PMDU1 ( // @[SIMDU.scala 454:21]
    .io_in_ready(PMDU1_io_in_ready),
    .io_in_valid(PMDU1_io_in_valid),
    .io_in_bits_DecodeIn_cf_pc(PMDU1_io_in_bits_DecodeIn_cf_pc),
    .io_in_bits_DecodeIn_cf_runahead_checkpoint_id(PMDU1_io_in_bits_DecodeIn_cf_runahead_checkpoint_id),
    .io_in_bits_DecodeIn_ctrl_fuOpType(PMDU1_io_in_bits_DecodeIn_ctrl_fuOpType),
    .io_in_bits_DecodeIn_ctrl_rfWen(PMDU1_io_in_bits_DecodeIn_ctrl_rfWen),
    .io_in_bits_DecodeIn_ctrl_rfDest(PMDU1_io_in_bits_DecodeIn_ctrl_rfDest),
    .io_in_bits_DecodeIn_data_src1(PMDU1_io_in_bits_DecodeIn_data_src1),
    .io_in_bits_DecodeIn_data_src2(PMDU1_io_in_bits_DecodeIn_data_src2),
    .io_in_bits_DecodeIn_data_src3(PMDU1_io_in_bits_DecodeIn_data_src3),
    .io_in_bits_DecodeIn_InstNo(PMDU1_io_in_bits_DecodeIn_InstNo),
    .io_in_bits_DecodeIn_InstFlag(PMDU1_io_in_bits_DecodeIn_InstFlag),
    .io_in_bits_Pctrl_isMul_16(PMDU1_io_in_bits_Pctrl_isMul_16),
    .io_in_bits_Pctrl_isMul_8(PMDU1_io_in_bits_Pctrl_isMul_8),
    .io_in_bits_Pctrl_isMSW_3232(PMDU1_io_in_bits_Pctrl_isMSW_3232),
    .io_in_bits_Pctrl_isMSW_3216(PMDU1_io_in_bits_Pctrl_isMSW_3216),
    .io_in_bits_Pctrl_isS1632(PMDU1_io_in_bits_Pctrl_isS1632),
    .io_in_bits_Pctrl_isS1664(PMDU1_io_in_bits_Pctrl_isS1664),
    .io_in_bits_Pctrl_is832(PMDU1_io_in_bits_Pctrl_is832),
    .io_in_bits_Pctrl_is3264(PMDU1_io_in_bits_Pctrl_is3264),
    .io_in_bits_Pctrl_is1664(PMDU1_io_in_bits_Pctrl_is1664),
    .io_in_bits_Pctrl_isQ15orQ31(PMDU1_io_in_bits_Pctrl_isQ15orQ31),
    .io_in_bits_Pctrl_isC31(PMDU1_io_in_bits_Pctrl_isC31),
    .io_in_bits_Pctrl_isQ15_64ONLY(PMDU1_io_in_bits_Pctrl_isQ15_64ONLY),
    .io_in_bits_Pctrl_isQ63_64ONLY(PMDU1_io_in_bits_Pctrl_isQ63_64ONLY),
    .io_in_bits_Pctrl_isMul_32_64ONLY(PMDU1_io_in_bits_Pctrl_isMul_32_64ONLY),
    .io_in_bits_Pctrl_isPMA_64ONLY(PMDU1_io_in_bits_Pctrl_isPMA_64ONLY),
    .io_in_bits_Pctrl_mulres9_0(PMDU1_io_in_bits_Pctrl_mulres9_0),
    .io_in_bits_Pctrl_mulres9_1(PMDU1_io_in_bits_Pctrl_mulres9_1),
    .io_in_bits_Pctrl_mulres9_2(PMDU1_io_in_bits_Pctrl_mulres9_2),
    .io_in_bits_Pctrl_mulres9_3(PMDU1_io_in_bits_Pctrl_mulres9_3),
    .io_in_bits_Pctrl_mulres17_0(PMDU1_io_in_bits_Pctrl_mulres17_0),
    .io_in_bits_Pctrl_mulres17_1(PMDU1_io_in_bits_Pctrl_mulres17_1),
    .io_in_bits_Pctrl_mulres33_0(PMDU1_io_in_bits_Pctrl_mulres33_0),
    .io_in_bits_Pctrl_mulres65_0(PMDU1_io_in_bits_Pctrl_mulres65_0),
    .io_out_ready(PMDU1_io_out_ready),
    .io_out_valid(PMDU1_io_out_valid),
    .io_out_bits_result(PMDU1_io_out_bits_result),
    .io_out_bits_DecodeOut_cf_pc(PMDU1_io_out_bits_DecodeOut_cf_pc),
    .io_out_bits_DecodeOut_cf_runahead_checkpoint_id(PMDU1_io_out_bits_DecodeOut_cf_runahead_checkpoint_id),
    .io_out_bits_DecodeOut_ctrl_fuOpType(PMDU1_io_out_bits_DecodeOut_ctrl_fuOpType),
    .io_out_bits_DecodeOut_ctrl_rfWen(PMDU1_io_out_bits_DecodeOut_ctrl_rfWen),
    .io_out_bits_DecodeOut_ctrl_rfDest(PMDU1_io_out_bits_DecodeOut_ctrl_rfDest),
    .io_out_bits_DecodeOut_data_src1(PMDU1_io_out_bits_DecodeOut_data_src1),
    .io_out_bits_DecodeOut_data_src2(PMDU1_io_out_bits_DecodeOut_data_src2),
    .io_out_bits_DecodeOut_data_src3(PMDU1_io_out_bits_DecodeOut_data_src3),
    .io_out_bits_DecodeOut_pext_OV(PMDU1_io_out_bits_DecodeOut_pext_OV),
    .io_out_bits_DecodeOut_InstNo(PMDU1_io_out_bits_DecodeOut_InstNo),
    .io_out_bits_DecodeOut_InstFlag(PMDU1_io_out_bits_DecodeOut_InstFlag),
    .io_FirstStageFire(PMDU1_io_FirstStageFire)
  );
  PIDU PIDU0 ( // @[SIMDU.scala 455:21]
    .io_DecodeIn_cf_instr(PIDU0_io_DecodeIn_cf_instr),
    .io_DecodeIn_cf_instrType(PIDU0_io_DecodeIn_cf_instrType),
    .io_DecodeIn_ctrl_fuOpType(PIDU0_io_DecodeIn_ctrl_fuOpType),
    .io_DecodeIn_ctrl_funct3(PIDU0_io_DecodeIn_ctrl_funct3),
    .io_DecodeIn_ctrl_func24(PIDU0_io_DecodeIn_ctrl_func24),
    .io_DecodeIn_ctrl_func23(PIDU0_io_DecodeIn_ctrl_func23),
    .io_DecodeIn_data_src1(PIDU0_io_DecodeIn_data_src1),
    .io_DecodeIn_data_src2(PIDU0_io_DecodeIn_data_src2),
    .io_Pctrl_isAdd_64(PIDU0_io_Pctrl_isAdd_64),
    .io_Pctrl_isAdd_32(PIDU0_io_Pctrl_isAdd_32),
    .io_Pctrl_isAdd_16(PIDU0_io_Pctrl_isAdd_16),
    .io_Pctrl_isAdd_8(PIDU0_io_Pctrl_isAdd_8),
    .io_Pctrl_isAdd_Q15(PIDU0_io_Pctrl_isAdd_Q15),
    .io_Pctrl_isAdd_Q31(PIDU0_io_Pctrl_isAdd_Q31),
    .io_Pctrl_isAdd_C31(PIDU0_io_Pctrl_isAdd_C31),
    .io_Pctrl_isAve(PIDU0_io_Pctrl_isAve),
    .io_Pctrl_isAdd(PIDU0_io_Pctrl_isAdd),
    .io_Pctrl_isSub_64(PIDU0_io_Pctrl_isSub_64),
    .io_Pctrl_isSub_32(PIDU0_io_Pctrl_isSub_32),
    .io_Pctrl_isSub_16(PIDU0_io_Pctrl_isSub_16),
    .io_Pctrl_isSub_8(PIDU0_io_Pctrl_isSub_8),
    .io_Pctrl_isSub_Q15(PIDU0_io_Pctrl_isSub_Q15),
    .io_Pctrl_isSub_Q31(PIDU0_io_Pctrl_isSub_Q31),
    .io_Pctrl_isSub_C31(PIDU0_io_Pctrl_isSub_C31),
    .io_Pctrl_isCras_16(PIDU0_io_Pctrl_isCras_16),
    .io_Pctrl_isCrsa_16(PIDU0_io_Pctrl_isCrsa_16),
    .io_Pctrl_isCras_32(PIDU0_io_Pctrl_isCras_32),
    .io_Pctrl_isCrsa_32(PIDU0_io_Pctrl_isCrsa_32),
    .io_Pctrl_isCr(PIDU0_io_Pctrl_isCr),
    .io_Pctrl_isStas_16(PIDU0_io_Pctrl_isStas_16),
    .io_Pctrl_isStsa_16(PIDU0_io_Pctrl_isStsa_16),
    .io_Pctrl_isStas_32(PIDU0_io_Pctrl_isStas_32),
    .io_Pctrl_isStsa_32(PIDU0_io_Pctrl_isStsa_32),
    .io_Pctrl_isSt(PIDU0_io_Pctrl_isSt),
    .io_Pctrl_isComp_16(PIDU0_io_Pctrl_isComp_16),
    .io_Pctrl_isComp_8(PIDU0_io_Pctrl_isComp_8),
    .io_Pctrl_isCompare(PIDU0_io_Pctrl_isCompare),
    .io_Pctrl_isMaxMin_16(PIDU0_io_Pctrl_isMaxMin_16),
    .io_Pctrl_isMaxMin_8(PIDU0_io_Pctrl_isMaxMin_8),
    .io_Pctrl_isMaxMin_XLEN(PIDU0_io_Pctrl_isMaxMin_XLEN),
    .io_Pctrl_isMaxMin_32(PIDU0_io_Pctrl_isMaxMin_32),
    .io_Pctrl_isMaxMin(PIDU0_io_Pctrl_isMaxMin),
    .io_Pctrl_isPbs(PIDU0_io_Pctrl_isPbs),
    .io_Pctrl_isRs_16(PIDU0_io_Pctrl_isRs_16),
    .io_Pctrl_isLs_16(PIDU0_io_Pctrl_isLs_16),
    .io_Pctrl_isLR_16(PIDU0_io_Pctrl_isLR_16),
    .io_Pctrl_isRs_8(PIDU0_io_Pctrl_isRs_8),
    .io_Pctrl_isLs_8(PIDU0_io_Pctrl_isLs_8),
    .io_Pctrl_isLR_8(PIDU0_io_Pctrl_isLR_8),
    .io_Pctrl_isRs_32(PIDU0_io_Pctrl_isRs_32),
    .io_Pctrl_isLs_32(PIDU0_io_Pctrl_isLs_32),
    .io_Pctrl_isLR_32(PIDU0_io_Pctrl_isLR_32),
    .io_Pctrl_isLR_Q31(PIDU0_io_Pctrl_isLR_Q31),
    .io_Pctrl_isLs_Q31(PIDU0_io_Pctrl_isLs_Q31),
    .io_Pctrl_isRs_XLEN(PIDU0_io_Pctrl_isRs_XLEN),
    .io_Pctrl_isSRAIWU(PIDU0_io_Pctrl_isSRAIWU),
    .io_Pctrl_isFSRW(PIDU0_io_Pctrl_isFSRW),
    .io_Pctrl_isWext(PIDU0_io_Pctrl_isWext),
    .io_Pctrl_isShifter(PIDU0_io_Pctrl_isShifter),
    .io_Pctrl_isClip_16(PIDU0_io_Pctrl_isClip_16),
    .io_Pctrl_isClip_8(PIDU0_io_Pctrl_isClip_8),
    .io_Pctrl_isclip_32(PIDU0_io_Pctrl_isclip_32),
    .io_Pctrl_isClip(PIDU0_io_Pctrl_isClip),
    .io_Pctrl_isSat_16(PIDU0_io_Pctrl_isSat_16),
    .io_Pctrl_isSat_8(PIDU0_io_Pctrl_isSat_8),
    .io_Pctrl_isSat_32(PIDU0_io_Pctrl_isSat_32),
    .io_Pctrl_isSat_W(PIDU0_io_Pctrl_isSat_W),
    .io_Pctrl_isSat(PIDU0_io_Pctrl_isSat),
    .io_Pctrl_isCnt_16(PIDU0_io_Pctrl_isCnt_16),
    .io_Pctrl_isCnt_8(PIDU0_io_Pctrl_isCnt_8),
    .io_Pctrl_isCnt_32(PIDU0_io_Pctrl_isCnt_32),
    .io_Pctrl_isCnt(PIDU0_io_Pctrl_isCnt),
    .io_Pctrl_isSwap_16(PIDU0_io_Pctrl_isSwap_16),
    .io_Pctrl_isSwap_8(PIDU0_io_Pctrl_isSwap_8),
    .io_Pctrl_isSwap(PIDU0_io_Pctrl_isSwap),
    .io_Pctrl_isUnpack(PIDU0_io_Pctrl_isUnpack),
    .io_Pctrl_isBitrev(PIDU0_io_Pctrl_isBitrev),
    .io_Pctrl_isCmix(PIDU0_io_Pctrl_isCmix),
    .io_Pctrl_isInsertb(PIDU0_io_Pctrl_isInsertb),
    .io_Pctrl_isPackbb(PIDU0_io_Pctrl_isPackbb),
    .io_Pctrl_isPackbt(PIDU0_io_Pctrl_isPackbt),
    .io_Pctrl_isPacktb(PIDU0_io_Pctrl_isPacktb),
    .io_Pctrl_isPacktt(PIDU0_io_Pctrl_isPacktt),
    .io_Pctrl_isPack(PIDU0_io_Pctrl_isPack),
    .io_Pctrl_isSub(PIDU0_io_Pctrl_isSub),
    .io_Pctrl_isAdder(PIDU0_io_Pctrl_isAdder),
    .io_Pctrl_SrcSigned(PIDU0_io_Pctrl_SrcSigned),
    .io_Pctrl_Saturating(PIDU0_io_Pctrl_Saturating),
    .io_Pctrl_Translation(PIDU0_io_Pctrl_Translation),
    .io_Pctrl_LessEqual(PIDU0_io_Pctrl_LessEqual),
    .io_Pctrl_LessThan(PIDU0_io_Pctrl_LessThan),
    .io_Pctrl_adderRes_ori(PIDU0_io_Pctrl_adderRes_ori),
    .io_Pctrl_adderRes(PIDU0_io_Pctrl_adderRes),
    .io_Pctrl_adderRes_ori_drophighestbit(PIDU0_io_Pctrl_adderRes_ori_drophighestbit),
    .io_Pctrl_Round(PIDU0_io_Pctrl_Round),
    .io_Pctrl_ShiftSigned(PIDU0_io_Pctrl_ShiftSigned),
    .io_Pctrl_Arithmetic(PIDU0_io_Pctrl_Arithmetic),
    .io_Pctrl_isMul_16(PIDU0_io_Pctrl_isMul_16),
    .io_Pctrl_isMul_8(PIDU0_io_Pctrl_isMul_8),
    .io_Pctrl_isMSW_3232(PIDU0_io_Pctrl_isMSW_3232),
    .io_Pctrl_isMSW_3216(PIDU0_io_Pctrl_isMSW_3216),
    .io_Pctrl_isS1632(PIDU0_io_Pctrl_isS1632),
    .io_Pctrl_isS1664(PIDU0_io_Pctrl_isS1664),
    .io_Pctrl_is832(PIDU0_io_Pctrl_is832),
    .io_Pctrl_is3264(PIDU0_io_Pctrl_is3264),
    .io_Pctrl_is1664(PIDU0_io_Pctrl_is1664),
    .io_Pctrl_isQ15orQ31(PIDU0_io_Pctrl_isQ15orQ31),
    .io_Pctrl_isC31(PIDU0_io_Pctrl_isC31),
    .io_Pctrl_isQ15_64ONLY(PIDU0_io_Pctrl_isQ15_64ONLY),
    .io_Pctrl_isQ63_64ONLY(PIDU0_io_Pctrl_isQ63_64ONLY),
    .io_Pctrl_isMul_32_64ONLY(PIDU0_io_Pctrl_isMul_32_64ONLY),
    .io_Pctrl_isPMA_64ONLY(PIDU0_io_Pctrl_isPMA_64ONLY),
    .io_Pctrl_mulres9_0(PIDU0_io_Pctrl_mulres9_0),
    .io_Pctrl_mulres9_1(PIDU0_io_Pctrl_mulres9_1),
    .io_Pctrl_mulres9_2(PIDU0_io_Pctrl_mulres9_2),
    .io_Pctrl_mulres9_3(PIDU0_io_Pctrl_mulres9_3),
    .io_Pctrl_mulres17_0(PIDU0_io_Pctrl_mulres17_0),
    .io_Pctrl_mulres17_1(PIDU0_io_Pctrl_mulres17_1),
    .io_Pctrl_mulres33_0(PIDU0_io_Pctrl_mulres33_0),
    .io_Pctrl_mulres65_0(PIDU0_io_Pctrl_mulres65_0)
  );
  PIDU_1 PIDU1 ( // @[SIMDU.scala 456:21]
    .io_DecodeIn_cf_instr(PIDU1_io_DecodeIn_cf_instr),
    .io_DecodeIn_cf_instrType(PIDU1_io_DecodeIn_cf_instrType),
    .io_DecodeIn_ctrl_fuOpType(PIDU1_io_DecodeIn_ctrl_fuOpType),
    .io_DecodeIn_ctrl_funct3(PIDU1_io_DecodeIn_ctrl_funct3),
    .io_DecodeIn_ctrl_func24(PIDU1_io_DecodeIn_ctrl_func24),
    .io_DecodeIn_ctrl_func23(PIDU1_io_DecodeIn_ctrl_func23),
    .io_DecodeIn_data_src1(PIDU1_io_DecodeIn_data_src1),
    .io_DecodeIn_data_src2(PIDU1_io_DecodeIn_data_src2),
    .io_Pctrl_isAdd_64(PIDU1_io_Pctrl_isAdd_64),
    .io_Pctrl_isAdd_32(PIDU1_io_Pctrl_isAdd_32),
    .io_Pctrl_isAdd_16(PIDU1_io_Pctrl_isAdd_16),
    .io_Pctrl_isAdd_8(PIDU1_io_Pctrl_isAdd_8),
    .io_Pctrl_isAdd_Q15(PIDU1_io_Pctrl_isAdd_Q15),
    .io_Pctrl_isAdd_Q31(PIDU1_io_Pctrl_isAdd_Q31),
    .io_Pctrl_isAdd_C31(PIDU1_io_Pctrl_isAdd_C31),
    .io_Pctrl_isAve(PIDU1_io_Pctrl_isAve),
    .io_Pctrl_isAdd(PIDU1_io_Pctrl_isAdd),
    .io_Pctrl_isSub_64(PIDU1_io_Pctrl_isSub_64),
    .io_Pctrl_isSub_32(PIDU1_io_Pctrl_isSub_32),
    .io_Pctrl_isSub_16(PIDU1_io_Pctrl_isSub_16),
    .io_Pctrl_isSub_8(PIDU1_io_Pctrl_isSub_8),
    .io_Pctrl_isSub_Q15(PIDU1_io_Pctrl_isSub_Q15),
    .io_Pctrl_isSub_Q31(PIDU1_io_Pctrl_isSub_Q31),
    .io_Pctrl_isSub_C31(PIDU1_io_Pctrl_isSub_C31),
    .io_Pctrl_isCras_16(PIDU1_io_Pctrl_isCras_16),
    .io_Pctrl_isCrsa_16(PIDU1_io_Pctrl_isCrsa_16),
    .io_Pctrl_isCras_32(PIDU1_io_Pctrl_isCras_32),
    .io_Pctrl_isCrsa_32(PIDU1_io_Pctrl_isCrsa_32),
    .io_Pctrl_isCr(PIDU1_io_Pctrl_isCr),
    .io_Pctrl_isStas_16(PIDU1_io_Pctrl_isStas_16),
    .io_Pctrl_isStsa_16(PIDU1_io_Pctrl_isStsa_16),
    .io_Pctrl_isStas_32(PIDU1_io_Pctrl_isStas_32),
    .io_Pctrl_isStsa_32(PIDU1_io_Pctrl_isStsa_32),
    .io_Pctrl_isSt(PIDU1_io_Pctrl_isSt),
    .io_Pctrl_isComp_16(PIDU1_io_Pctrl_isComp_16),
    .io_Pctrl_isComp_8(PIDU1_io_Pctrl_isComp_8),
    .io_Pctrl_isCompare(PIDU1_io_Pctrl_isCompare),
    .io_Pctrl_isMaxMin_16(PIDU1_io_Pctrl_isMaxMin_16),
    .io_Pctrl_isMaxMin_8(PIDU1_io_Pctrl_isMaxMin_8),
    .io_Pctrl_isMaxMin_XLEN(PIDU1_io_Pctrl_isMaxMin_XLEN),
    .io_Pctrl_isMaxMin_32(PIDU1_io_Pctrl_isMaxMin_32),
    .io_Pctrl_isMaxMin(PIDU1_io_Pctrl_isMaxMin),
    .io_Pctrl_isPbs(PIDU1_io_Pctrl_isPbs),
    .io_Pctrl_isRs_16(PIDU1_io_Pctrl_isRs_16),
    .io_Pctrl_isLs_16(PIDU1_io_Pctrl_isLs_16),
    .io_Pctrl_isLR_16(PIDU1_io_Pctrl_isLR_16),
    .io_Pctrl_isRs_8(PIDU1_io_Pctrl_isRs_8),
    .io_Pctrl_isLs_8(PIDU1_io_Pctrl_isLs_8),
    .io_Pctrl_isLR_8(PIDU1_io_Pctrl_isLR_8),
    .io_Pctrl_isRs_32(PIDU1_io_Pctrl_isRs_32),
    .io_Pctrl_isLs_32(PIDU1_io_Pctrl_isLs_32),
    .io_Pctrl_isLR_32(PIDU1_io_Pctrl_isLR_32),
    .io_Pctrl_isLR_Q31(PIDU1_io_Pctrl_isLR_Q31),
    .io_Pctrl_isLs_Q31(PIDU1_io_Pctrl_isLs_Q31),
    .io_Pctrl_isRs_XLEN(PIDU1_io_Pctrl_isRs_XLEN),
    .io_Pctrl_isSRAIWU(PIDU1_io_Pctrl_isSRAIWU),
    .io_Pctrl_isFSRW(PIDU1_io_Pctrl_isFSRW),
    .io_Pctrl_isWext(PIDU1_io_Pctrl_isWext),
    .io_Pctrl_isShifter(PIDU1_io_Pctrl_isShifter),
    .io_Pctrl_isClip_16(PIDU1_io_Pctrl_isClip_16),
    .io_Pctrl_isClip_8(PIDU1_io_Pctrl_isClip_8),
    .io_Pctrl_isclip_32(PIDU1_io_Pctrl_isclip_32),
    .io_Pctrl_isClip(PIDU1_io_Pctrl_isClip),
    .io_Pctrl_isSat_16(PIDU1_io_Pctrl_isSat_16),
    .io_Pctrl_isSat_8(PIDU1_io_Pctrl_isSat_8),
    .io_Pctrl_isSat_32(PIDU1_io_Pctrl_isSat_32),
    .io_Pctrl_isSat_W(PIDU1_io_Pctrl_isSat_W),
    .io_Pctrl_isSat(PIDU1_io_Pctrl_isSat),
    .io_Pctrl_isCnt_16(PIDU1_io_Pctrl_isCnt_16),
    .io_Pctrl_isCnt_8(PIDU1_io_Pctrl_isCnt_8),
    .io_Pctrl_isCnt_32(PIDU1_io_Pctrl_isCnt_32),
    .io_Pctrl_isCnt(PIDU1_io_Pctrl_isCnt),
    .io_Pctrl_isSwap_16(PIDU1_io_Pctrl_isSwap_16),
    .io_Pctrl_isSwap_8(PIDU1_io_Pctrl_isSwap_8),
    .io_Pctrl_isSwap(PIDU1_io_Pctrl_isSwap),
    .io_Pctrl_isUnpack(PIDU1_io_Pctrl_isUnpack),
    .io_Pctrl_isBitrev(PIDU1_io_Pctrl_isBitrev),
    .io_Pctrl_isCmix(PIDU1_io_Pctrl_isCmix),
    .io_Pctrl_isInsertb(PIDU1_io_Pctrl_isInsertb),
    .io_Pctrl_isPackbb(PIDU1_io_Pctrl_isPackbb),
    .io_Pctrl_isPackbt(PIDU1_io_Pctrl_isPackbt),
    .io_Pctrl_isPacktb(PIDU1_io_Pctrl_isPacktb),
    .io_Pctrl_isPacktt(PIDU1_io_Pctrl_isPacktt),
    .io_Pctrl_isPack(PIDU1_io_Pctrl_isPack),
    .io_Pctrl_isSub(PIDU1_io_Pctrl_isSub),
    .io_Pctrl_isAdder(PIDU1_io_Pctrl_isAdder),
    .io_Pctrl_SrcSigned(PIDU1_io_Pctrl_SrcSigned),
    .io_Pctrl_Saturating(PIDU1_io_Pctrl_Saturating),
    .io_Pctrl_Translation(PIDU1_io_Pctrl_Translation),
    .io_Pctrl_LessEqual(PIDU1_io_Pctrl_LessEqual),
    .io_Pctrl_LessThan(PIDU1_io_Pctrl_LessThan),
    .io_Pctrl_adderRes_ori(PIDU1_io_Pctrl_adderRes_ori),
    .io_Pctrl_adderRes(PIDU1_io_Pctrl_adderRes),
    .io_Pctrl_adderRes_ori_drophighestbit(PIDU1_io_Pctrl_adderRes_ori_drophighestbit),
    .io_Pctrl_Round(PIDU1_io_Pctrl_Round),
    .io_Pctrl_ShiftSigned(PIDU1_io_Pctrl_ShiftSigned),
    .io_Pctrl_Arithmetic(PIDU1_io_Pctrl_Arithmetic),
    .io_Pctrl_isMul_16(PIDU1_io_Pctrl_isMul_16),
    .io_Pctrl_isMul_8(PIDU1_io_Pctrl_isMul_8),
    .io_Pctrl_isMSW_3232(PIDU1_io_Pctrl_isMSW_3232),
    .io_Pctrl_isMSW_3216(PIDU1_io_Pctrl_isMSW_3216),
    .io_Pctrl_isS1632(PIDU1_io_Pctrl_isS1632),
    .io_Pctrl_isS1664(PIDU1_io_Pctrl_isS1664),
    .io_Pctrl_is832(PIDU1_io_Pctrl_is832),
    .io_Pctrl_is3264(PIDU1_io_Pctrl_is3264),
    .io_Pctrl_is1664(PIDU1_io_Pctrl_is1664),
    .io_Pctrl_isQ15orQ31(PIDU1_io_Pctrl_isQ15orQ31),
    .io_Pctrl_isC31(PIDU1_io_Pctrl_isC31),
    .io_Pctrl_isQ15_64ONLY(PIDU1_io_Pctrl_isQ15_64ONLY),
    .io_Pctrl_isQ63_64ONLY(PIDU1_io_Pctrl_isQ63_64ONLY),
    .io_Pctrl_isMul_32_64ONLY(PIDU1_io_Pctrl_isMul_32_64ONLY),
    .io_Pctrl_isPMA_64ONLY(PIDU1_io_Pctrl_isPMA_64ONLY),
    .io_Pctrl_mulres9_0(PIDU1_io_Pctrl_mulres9_0),
    .io_Pctrl_mulres9_1(PIDU1_io_Pctrl_mulres9_1),
    .io_Pctrl_mulres9_2(PIDU1_io_Pctrl_mulres9_2),
    .io_Pctrl_mulres9_3(PIDU1_io_Pctrl_mulres9_3),
    .io_Pctrl_mulres17_0(PIDU1_io_Pctrl_mulres17_0),
    .io_Pctrl_mulres17_1(PIDU1_io_Pctrl_mulres17_1),
    .io_Pctrl_mulres33_0(PIDU1_io_Pctrl_mulres33_0),
    .io_Pctrl_mulres65_0(PIDU1_io_Pctrl_mulres65_0)
  );
  assign io_DecodeOut_0_cf_pc = _T_95 ? PALU0_io_out_bits_DecodeOut_cf_pc : _GEN_4759; // @[SIMDU.scala 617:21 619:20]
  assign io_DecodeOut_0_cf_runahead_checkpoint_id = _T_95 ? PALU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id :
    _GEN_4723; // @[SIMDU.scala 617:21 619:20]
  assign io_DecodeOut_0_ctrl_rfWen = _T_95 ? PALU0_io_out_bits_DecodeOut_ctrl_rfWen : _GEN_4710; // @[SIMDU.scala 617:21 619:20]
  assign io_DecodeOut_0_ctrl_rfDest = _T_95 ? PALU0_io_out_bits_DecodeOut_ctrl_rfDest : _GEN_4709; // @[SIMDU.scala 617:21 619:20]
  assign io_DecodeOut_0_pext_OV = _T_95 ? PALU0_io_out_bits_DecodeOut_pext_OV : _GEN_4697; // @[SIMDU.scala 617:21 619:20]
  assign io_DecodeOut_0_InstNo = _T_95 ? PALU0_io_out_bits_DecodeOut_InstNo : _GEN_4696; // @[SIMDU.scala 617:21 619:20]
  assign io_DecodeOut_1_cf_pc = queen == 2'h0 ? PALU0_io_out_bits_DecodeOut_cf_pc : _GEN_4972; // @[SIMDU.scala 638:22 640:20]
  assign io_DecodeOut_1_cf_runahead_checkpoint_id = queen == 2'h0 ?
    PALU0_io_out_bits_DecodeOut_cf_runahead_checkpoint_id : _GEN_4936; // @[SIMDU.scala 638:22 640:20]
  assign io_DecodeOut_1_ctrl_rfWen = queen == 2'h0 ? PALU0_io_out_bits_DecodeOut_ctrl_rfWen : _GEN_4923; // @[SIMDU.scala 638:22 640:20]
  assign io_DecodeOut_1_ctrl_rfDest = queen == 2'h0 ? PALU0_io_out_bits_DecodeOut_ctrl_rfDest : _GEN_4922; // @[SIMDU.scala 638:22 640:20]
  assign io_DecodeOut_1_pext_OV = queen == 2'h0 ? PALU0_io_out_bits_DecodeOut_pext_OV : _GEN_4910; // @[SIMDU.scala 638:22 640:20]
  assign io_DecodeOut_1_InstNo = queen == 2'h0 ? PALU0_io_out_bits_DecodeOut_InstNo : _GEN_4909; // @[SIMDU.scala 638:22 640:20]
  assign io_FirstStageFire_0 = _GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15) ? _GEN_2816 :
    _GEN_3721; // @[SIMDU.scala 547:184]
  assign io_FirstStageFire_1 = _GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15) ? _GEN_2817 :
    _GEN_3722; // @[SIMDU.scala 547:184]
  assign io_in_0_ready = ~io_in_0_valid | io_FirstStageFire_0; // @[SIMDU.scala 458:29]
  assign io_in_1_ready = ~io_in_1_valid | io_FirstStageFire_1; // @[SIMDU.scala 459:29]
  assign io_out_0_valid = _T_95 ? PALU0_io_out_valid : _GEN_4761; // @[SIMDU.scala 617:21 620:20]
  assign io_out_0_bits = _T_95 ? PALU0_io_out_bits_result : _GEN_4694; // @[SIMDU.scala 617:21 618:20]
  assign io_out_1_valid = queen == 2'h0 ? PALU0_io_out_valid : _GEN_4974; // @[SIMDU.scala 638:22 641:20]
  assign io_out_1_bits = queen == 2'h0 ? PALU0_io_out_bits_result : _GEN_4907; // @[SIMDU.scala 638:22 639:20]
  assign PALU0_io_in_valid = PALU0_valid; // @[SIMDU.scala 575:21]
  assign PALU0_io_in_bits_DecodeIn_cf_pc = PALU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_cf_runahead_checkpoint_id = PALU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_ctrl_fuOpType = PALU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_ctrl_funct3 = PALU0_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_ctrl_func24 = PALU0_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_ctrl_rfWen = PALU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_ctrl_rfDest = PALU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_data_src1 = PALU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_data_src2 = PALU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_data_src3 = PALU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_InstNo = PALU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_DecodeIn_InstFlag = PALU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_64 = PALU0_bits_Pctrl_isAdd_64; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_32 = PALU0_bits_Pctrl_isAdd_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_16 = PALU0_bits_Pctrl_isAdd_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_8 = PALU0_bits_Pctrl_isAdd_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_Q15 = PALU0_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_Q31 = PALU0_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdd_C31 = PALU0_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAve = PALU0_bits_Pctrl_isAve; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_64 = PALU0_bits_Pctrl_isSub_64; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_32 = PALU0_bits_Pctrl_isSub_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_16 = PALU0_bits_Pctrl_isSub_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_8 = PALU0_bits_Pctrl_isSub_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_Q15 = PALU0_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_Q31 = PALU0_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub_C31 = PALU0_bits_Pctrl_isSub_C31; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCras_16 = PALU0_bits_Pctrl_isCras_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCrsa_16 = PALU0_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCras_32 = PALU0_bits_Pctrl_isCras_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCrsa_32 = PALU0_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isStas_16 = PALU0_bits_Pctrl_isStas_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isStsa_16 = PALU0_bits_Pctrl_isStsa_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isStas_32 = PALU0_bits_Pctrl_isStas_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isStsa_32 = PALU0_bits_Pctrl_isStsa_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isComp_16 = PALU0_bits_Pctrl_isComp_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isComp_8 = PALU0_bits_Pctrl_isComp_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCompare = PALU0_bits_Pctrl_isCompare; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isMaxMin_16 = PALU0_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isMaxMin_8 = PALU0_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isMaxMin_XLEN = PALU0_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isMaxMin_32 = PALU0_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isMaxMin = PALU0_bits_Pctrl_isMaxMin; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isPbs = PALU0_bits_Pctrl_isPbs; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isRs_16 = PALU0_bits_Pctrl_isRs_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLs_16 = PALU0_bits_Pctrl_isLs_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLR_16 = PALU0_bits_Pctrl_isLR_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isRs_8 = PALU0_bits_Pctrl_isRs_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLs_8 = PALU0_bits_Pctrl_isLs_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLR_8 = PALU0_bits_Pctrl_isLR_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isRs_32 = PALU0_bits_Pctrl_isRs_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLs_32 = PALU0_bits_Pctrl_isLs_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLR_32 = PALU0_bits_Pctrl_isLR_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLR_Q31 = PALU0_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isLs_Q31 = PALU0_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isRs_XLEN = PALU0_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSRAIWU = PALU0_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isFSRW = PALU0_bits_Pctrl_isFSRW; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isWext = PALU0_bits_Pctrl_isWext; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isShifter = PALU0_bits_Pctrl_isShifter; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isClip_16 = PALU0_bits_Pctrl_isClip_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isClip_8 = PALU0_bits_Pctrl_isClip_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isclip_32 = PALU0_bits_Pctrl_isclip_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isClip = PALU0_bits_Pctrl_isClip; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSat_16 = PALU0_bits_Pctrl_isSat_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSat_8 = PALU0_bits_Pctrl_isSat_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSat_32 = PALU0_bits_Pctrl_isSat_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSat_W = PALU0_bits_Pctrl_isSat_W; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSat = PALU0_bits_Pctrl_isSat; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCnt_16 = PALU0_bits_Pctrl_isCnt_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCnt_8 = PALU0_bits_Pctrl_isCnt_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCnt_32 = PALU0_bits_Pctrl_isCnt_32; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCnt = PALU0_bits_Pctrl_isCnt; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSwap_16 = PALU0_bits_Pctrl_isSwap_16; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSwap_8 = PALU0_bits_Pctrl_isSwap_8; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSwap = PALU0_bits_Pctrl_isSwap; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isUnpack = PALU0_bits_Pctrl_isUnpack; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isBitrev = PALU0_bits_Pctrl_isBitrev; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isCmix = PALU0_bits_Pctrl_isCmix; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isInsertb = PALU0_bits_Pctrl_isInsertb; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isPackbb = PALU0_bits_Pctrl_isPackbb; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isPackbt = PALU0_bits_Pctrl_isPackbt; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isPacktb = PALU0_bits_Pctrl_isPacktb; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isPacktt = PALU0_bits_Pctrl_isPacktt; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isPack = PALU0_bits_Pctrl_isPack; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isSub = PALU0_bits_Pctrl_isSub; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_isAdder = PALU0_bits_Pctrl_isAdder; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_SrcSigned = PALU0_bits_Pctrl_SrcSigned; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_Saturating = PALU0_bits_Pctrl_Saturating; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_Translation = PALU0_bits_Pctrl_Translation; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_LessEqual = PALU0_bits_Pctrl_LessEqual; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_LessThan = PALU0_bits_Pctrl_LessThan; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_adderRes_ori = PALU0_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_adderRes = PALU0_bits_Pctrl_adderRes; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_adderRes_ori_drophighestbit = PALU0_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_Round = PALU0_bits_Pctrl_Round; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_ShiftSigned = PALU0_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 576:21]
  assign PALU0_io_in_bits_Pctrl_Arithmetic = PALU0_bits_Pctrl_Arithmetic; // @[SIMDU.scala 576:21]
  assign PALU0_io_out_ready = queen == 2'h0 ? io_out_1_ready : _GEN_4833; // @[SIMDU.scala 638:22 642:24]
  assign PMDU0_io_in_valid = PMDU0_valid; // @[SIMDU.scala 585:21]
  assign PMDU0_io_in_bits_DecodeIn_cf_pc = PMDU0_bits_DecodeIn_cf_pc; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_cf_runahead_checkpoint_id = PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_ctrl_fuOpType = PMDU0_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_ctrl_rfWen = PMDU0_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_ctrl_rfDest = PMDU0_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_data_src1 = PMDU0_bits_DecodeIn_data_src1; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_data_src2 = PMDU0_bits_DecodeIn_data_src2; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_data_src3 = PMDU0_bits_DecodeIn_data_src3; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_InstNo = PMDU0_bits_DecodeIn_InstNo; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_DecodeIn_InstFlag = PMDU0_bits_DecodeIn_InstFlag; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isMul_16 = PMDU0_bits_Pctrl_isMul_16; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isMul_8 = PMDU0_bits_Pctrl_isMul_8; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isMSW_3232 = PMDU0_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isMSW_3216 = PMDU0_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isS1632 = PMDU0_bits_Pctrl_isS1632; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isS1664 = PMDU0_bits_Pctrl_isS1664; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_is832 = PMDU0_bits_Pctrl_is832; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_is3264 = PMDU0_bits_Pctrl_is3264; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_is1664 = PMDU0_bits_Pctrl_is1664; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isQ15orQ31 = PMDU0_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isC31 = PMDU0_bits_Pctrl_isC31; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isQ15_64ONLY = PMDU0_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isQ63_64ONLY = PMDU0_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isMul_32_64ONLY = PMDU0_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_isPMA_64ONLY = PMDU0_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres9_0 = PMDU0_bits_Pctrl_mulres9_0; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres9_1 = PMDU0_bits_Pctrl_mulres9_1; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres9_2 = PMDU0_bits_Pctrl_mulres9_2; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres9_3 = PMDU0_bits_Pctrl_mulres9_3; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres17_0 = PMDU0_bits_Pctrl_mulres17_0; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres17_1 = PMDU0_bits_Pctrl_mulres17_1; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres33_0 = PMDU0_bits_Pctrl_mulres33_0; // @[SIMDU.scala 586:21]
  assign PMDU0_io_in_bits_Pctrl_mulres65_0 = PMDU0_bits_Pctrl_mulres65_0; // @[SIMDU.scala 586:21]
  assign PMDU0_io_out_ready = queen == 2'h0 ? _GEN_4835 : _GEN_4976; // @[SIMDU.scala 638:22]
  assign PALU1_io_in_valid = PALU1_valid; // @[SIMDU.scala 580:21]
  assign PALU1_io_in_bits_DecodeIn_cf_pc = PALU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_cf_runahead_checkpoint_id = PALU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_ctrl_fuOpType = PALU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_ctrl_funct3 = PALU1_bits_DecodeIn_ctrl_funct3; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_ctrl_func24 = PALU1_bits_DecodeIn_ctrl_func24; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_ctrl_rfWen = PALU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_ctrl_rfDest = PALU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_data_src1 = PALU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_data_src2 = PALU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_data_src3 = PALU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_InstNo = PALU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_DecodeIn_InstFlag = PALU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_64 = PALU1_bits_Pctrl_isAdd_64; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_32 = PALU1_bits_Pctrl_isAdd_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_16 = PALU1_bits_Pctrl_isAdd_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_8 = PALU1_bits_Pctrl_isAdd_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_Q15 = PALU1_bits_Pctrl_isAdd_Q15; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_Q31 = PALU1_bits_Pctrl_isAdd_Q31; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdd_C31 = PALU1_bits_Pctrl_isAdd_C31; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAve = PALU1_bits_Pctrl_isAve; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_64 = PALU1_bits_Pctrl_isSub_64; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_32 = PALU1_bits_Pctrl_isSub_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_16 = PALU1_bits_Pctrl_isSub_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_8 = PALU1_bits_Pctrl_isSub_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_Q15 = PALU1_bits_Pctrl_isSub_Q15; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_Q31 = PALU1_bits_Pctrl_isSub_Q31; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub_C31 = PALU1_bits_Pctrl_isSub_C31; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCras_16 = PALU1_bits_Pctrl_isCras_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCrsa_16 = PALU1_bits_Pctrl_isCrsa_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCras_32 = PALU1_bits_Pctrl_isCras_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCrsa_32 = PALU1_bits_Pctrl_isCrsa_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isStas_16 = PALU1_bits_Pctrl_isStas_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isStsa_16 = PALU1_bits_Pctrl_isStsa_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isStas_32 = PALU1_bits_Pctrl_isStas_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isStsa_32 = PALU1_bits_Pctrl_isStsa_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isComp_16 = PALU1_bits_Pctrl_isComp_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isComp_8 = PALU1_bits_Pctrl_isComp_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCompare = PALU1_bits_Pctrl_isCompare; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isMaxMin_16 = PALU1_bits_Pctrl_isMaxMin_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isMaxMin_8 = PALU1_bits_Pctrl_isMaxMin_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isMaxMin_XLEN = PALU1_bits_Pctrl_isMaxMin_XLEN; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isMaxMin_32 = PALU1_bits_Pctrl_isMaxMin_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isMaxMin = PALU1_bits_Pctrl_isMaxMin; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isPbs = PALU1_bits_Pctrl_isPbs; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isRs_16 = PALU1_bits_Pctrl_isRs_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLs_16 = PALU1_bits_Pctrl_isLs_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLR_16 = PALU1_bits_Pctrl_isLR_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isRs_8 = PALU1_bits_Pctrl_isRs_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLs_8 = PALU1_bits_Pctrl_isLs_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLR_8 = PALU1_bits_Pctrl_isLR_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isRs_32 = PALU1_bits_Pctrl_isRs_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLs_32 = PALU1_bits_Pctrl_isLs_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLR_32 = PALU1_bits_Pctrl_isLR_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLR_Q31 = PALU1_bits_Pctrl_isLR_Q31; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isLs_Q31 = PALU1_bits_Pctrl_isLs_Q31; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isRs_XLEN = PALU1_bits_Pctrl_isRs_XLEN; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSRAIWU = PALU1_bits_Pctrl_isSRAIWU; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isFSRW = PALU1_bits_Pctrl_isFSRW; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isWext = PALU1_bits_Pctrl_isWext; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isShifter = PALU1_bits_Pctrl_isShifter; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isClip_16 = PALU1_bits_Pctrl_isClip_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isClip_8 = PALU1_bits_Pctrl_isClip_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isclip_32 = PALU1_bits_Pctrl_isclip_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isClip = PALU1_bits_Pctrl_isClip; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSat_16 = PALU1_bits_Pctrl_isSat_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSat_8 = PALU1_bits_Pctrl_isSat_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSat_32 = PALU1_bits_Pctrl_isSat_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSat_W = PALU1_bits_Pctrl_isSat_W; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSat = PALU1_bits_Pctrl_isSat; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCnt_16 = PALU1_bits_Pctrl_isCnt_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCnt_8 = PALU1_bits_Pctrl_isCnt_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCnt_32 = PALU1_bits_Pctrl_isCnt_32; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCnt = PALU1_bits_Pctrl_isCnt; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSwap_16 = PALU1_bits_Pctrl_isSwap_16; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSwap_8 = PALU1_bits_Pctrl_isSwap_8; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSwap = PALU1_bits_Pctrl_isSwap; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isUnpack = PALU1_bits_Pctrl_isUnpack; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isBitrev = PALU1_bits_Pctrl_isBitrev; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isCmix = PALU1_bits_Pctrl_isCmix; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isInsertb = PALU1_bits_Pctrl_isInsertb; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isPackbb = PALU1_bits_Pctrl_isPackbb; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isPackbt = PALU1_bits_Pctrl_isPackbt; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isPacktb = PALU1_bits_Pctrl_isPacktb; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isPacktt = PALU1_bits_Pctrl_isPacktt; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isPack = PALU1_bits_Pctrl_isPack; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isSub = PALU1_bits_Pctrl_isSub; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_isAdder = PALU1_bits_Pctrl_isAdder; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_SrcSigned = PALU1_bits_Pctrl_SrcSigned; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_Saturating = PALU1_bits_Pctrl_Saturating; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_Translation = PALU1_bits_Pctrl_Translation; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_LessEqual = PALU1_bits_Pctrl_LessEqual; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_LessThan = PALU1_bits_Pctrl_LessThan; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_adderRes_ori = PALU1_bits_Pctrl_adderRes_ori; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_adderRes = PALU1_bits_Pctrl_adderRes; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_adderRes_ori_drophighestbit = PALU1_bits_Pctrl_adderRes_ori_drophighestbit; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_Round = PALU1_bits_Pctrl_Round; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_ShiftSigned = PALU1_bits_Pctrl_ShiftSigned; // @[SIMDU.scala 581:21]
  assign PALU1_io_in_bits_Pctrl_Arithmetic = PALU1_bits_Pctrl_Arithmetic; // @[SIMDU.scala 581:21]
  assign PALU1_io_out_ready = queen == 2'h0 ? _GEN_4834 : _GEN_4975; // @[SIMDU.scala 638:22]
  assign PMDU1_io_in_valid = PMDU1_valid; // @[SIMDU.scala 591:21]
  assign PMDU1_io_in_bits_DecodeIn_cf_pc = PMDU1_bits_DecodeIn_cf_pc; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_cf_runahead_checkpoint_id = PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_ctrl_fuOpType = PMDU1_bits_DecodeIn_ctrl_fuOpType; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_ctrl_rfWen = PMDU1_bits_DecodeIn_ctrl_rfWen; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_ctrl_rfDest = PMDU1_bits_DecodeIn_ctrl_rfDest; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_data_src1 = PMDU1_bits_DecodeIn_data_src1; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_data_src2 = PMDU1_bits_DecodeIn_data_src2; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_data_src3 = PMDU1_bits_DecodeIn_data_src3; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_InstNo = PMDU1_bits_DecodeIn_InstNo; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_DecodeIn_InstFlag = PMDU1_bits_DecodeIn_InstFlag; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isMul_16 = PMDU1_bits_Pctrl_isMul_16; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isMul_8 = PMDU1_bits_Pctrl_isMul_8; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isMSW_3232 = PMDU1_bits_Pctrl_isMSW_3232; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isMSW_3216 = PMDU1_bits_Pctrl_isMSW_3216; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isS1632 = PMDU1_bits_Pctrl_isS1632; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isS1664 = PMDU1_bits_Pctrl_isS1664; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_is832 = PMDU1_bits_Pctrl_is832; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_is3264 = PMDU1_bits_Pctrl_is3264; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_is1664 = PMDU1_bits_Pctrl_is1664; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isQ15orQ31 = PMDU1_bits_Pctrl_isQ15orQ31; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isC31 = PMDU1_bits_Pctrl_isC31; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isQ15_64ONLY = PMDU1_bits_Pctrl_isQ15_64ONLY; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isQ63_64ONLY = PMDU1_bits_Pctrl_isQ63_64ONLY; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isMul_32_64ONLY = PMDU1_bits_Pctrl_isMul_32_64ONLY; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_isPMA_64ONLY = PMDU1_bits_Pctrl_isPMA_64ONLY; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres9_0 = PMDU1_bits_Pctrl_mulres9_0; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres9_1 = PMDU1_bits_Pctrl_mulres9_1; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres9_2 = PMDU1_bits_Pctrl_mulres9_2; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres9_3 = PMDU1_bits_Pctrl_mulres9_3; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres17_0 = PMDU1_bits_Pctrl_mulres17_0; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres17_1 = PMDU1_bits_Pctrl_mulres17_1; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres33_0 = PMDU1_bits_Pctrl_mulres33_0; // @[SIMDU.scala 592:21]
  assign PMDU1_io_in_bits_Pctrl_mulres65_0 = PMDU1_bits_Pctrl_mulres65_0; // @[SIMDU.scala 592:21]
  assign PMDU1_io_out_ready = queen == 2'h0 ? _GEN_4836 : _GEN_4977; // @[SIMDU.scala 638:22]
  assign PIDU0_io_DecodeIn_cf_instr = io_DecodeIn_0_cf_instr; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_cf_instrType = io_DecodeIn_0_cf_instrType; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_ctrl_fuOpType = io_DecodeIn_0_ctrl_fuOpType; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_ctrl_funct3 = io_DecodeIn_0_ctrl_funct3; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_ctrl_func24 = io_DecodeIn_0_ctrl_func24; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_ctrl_func23 = io_DecodeIn_0_ctrl_func23; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_data_src1 = io_DecodeIn_0_data_src1; // @[SIMDU.scala 477:21]
  assign PIDU0_io_DecodeIn_data_src2 = io_DecodeIn_0_data_src2; // @[SIMDU.scala 477:21]
  assign PIDU1_io_DecodeIn_cf_instr = io_DecodeIn_1_cf_instr; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_cf_instrType = io_DecodeIn_1_cf_instrType; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_ctrl_fuOpType = io_DecodeIn_1_ctrl_fuOpType; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_ctrl_funct3 = io_DecodeIn_1_ctrl_funct3; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_ctrl_func24 = io_DecodeIn_1_ctrl_func24; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_ctrl_func23 = io_DecodeIn_1_ctrl_func23; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_data_src1 = io_DecodeIn_1_data_src1; // @[SIMDU.scala 478:21]
  assign PIDU1_io_DecodeIn_data_src2 = io_DecodeIn_1_data_src2; // @[SIMDU.scala 478:21]
  always @(posedge clock) begin
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_cf_pc <= 39'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_cf_pc <= io_DecodeIn_1_cf_pc; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_cf_pc <= io_DecodeIn_0_cf_pc;
        end
      end else begin
        PALU0_bits_DecodeIn_cf_pc <= _GEN_1662;
      end
    end else begin
      PALU0_bits_DecodeIn_cf_pc <= _GEN_1662;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_cf_runahead_checkpoint_id <= 64'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_cf_runahead_checkpoint_id <= io_DecodeIn_1_cf_runahead_checkpoint_id; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_cf_runahead_checkpoint_id <= io_DecodeIn_0_cf_runahead_checkpoint_id;
        end
      end else begin
        PALU0_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1626;
      end
    end else begin
      PALU0_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1626;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_ctrl_fuOpType <= 7'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_ctrl_fuOpType <= io_DecodeIn_1_ctrl_fuOpType; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_ctrl_fuOpType <= io_DecodeIn_0_ctrl_fuOpType;
        end
      end else begin
        PALU0_bits_DecodeIn_ctrl_fuOpType <= _GEN_1620;
      end
    end else begin
      PALU0_bits_DecodeIn_ctrl_fuOpType <= _GEN_1620;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_ctrl_funct3 <= 3'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_ctrl_funct3 <= io_DecodeIn_1_ctrl_funct3; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_ctrl_funct3 <= io_DecodeIn_0_ctrl_funct3;
        end
      end else begin
        PALU0_bits_DecodeIn_ctrl_funct3 <= _GEN_1619;
      end
    end else begin
      PALU0_bits_DecodeIn_ctrl_funct3 <= _GEN_1619;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_ctrl_func24 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_ctrl_func24 <= io_DecodeIn_1_ctrl_func24; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_ctrl_func24 <= io_DecodeIn_0_ctrl_func24;
        end
      end else begin
        PALU0_bits_DecodeIn_ctrl_func24 <= _GEN_1618;
      end
    end else begin
      PALU0_bits_DecodeIn_ctrl_func24 <= _GEN_1618;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_ctrl_rfWen <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_ctrl_rfWen <= io_DecodeIn_1_ctrl_rfWen; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_ctrl_rfWen <= io_DecodeIn_0_ctrl_rfWen;
        end
      end else begin
        PALU0_bits_DecodeIn_ctrl_rfWen <= _GEN_1613;
      end
    end else begin
      PALU0_bits_DecodeIn_ctrl_rfWen <= _GEN_1613;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_ctrl_rfDest <= 5'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_ctrl_rfDest <= io_DecodeIn_1_ctrl_rfDest; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_ctrl_rfDest <= io_DecodeIn_0_ctrl_rfDest;
        end
      end else begin
        PALU0_bits_DecodeIn_ctrl_rfDest <= _GEN_1612;
      end
    end else begin
      PALU0_bits_DecodeIn_ctrl_rfDest <= _GEN_1612;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_data_src1 <= 64'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_data_src1 <= io_DecodeIn_1_data_src1; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_data_src1 <= io_DecodeIn_0_data_src1;
        end
      end else begin
        PALU0_bits_DecodeIn_data_src1 <= _GEN_1604;
      end
    end else begin
      PALU0_bits_DecodeIn_data_src1 <= _GEN_1604;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_data_src2 <= 64'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_data_src2 <= io_DecodeIn_1_data_src2; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_data_src2 <= io_DecodeIn_0_data_src2;
        end
      end else begin
        PALU0_bits_DecodeIn_data_src2 <= _GEN_1603;
      end
    end else begin
      PALU0_bits_DecodeIn_data_src2 <= _GEN_1603;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_data_src3 <= 64'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_data_src3 <= io_DecodeIn_1_data_src3; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_data_src3 <= io_DecodeIn_0_data_src3;
        end
      end else begin
        PALU0_bits_DecodeIn_data_src3 <= _GEN_1602;
      end
    end else begin
      PALU0_bits_DecodeIn_data_src3 <= _GEN_1602;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_InstNo <= 5'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_InstNo <= io_DecodeIn_1_InstNo; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_InstNo <= io_DecodeIn_0_InstNo;
        end
      end else begin
        PALU0_bits_DecodeIn_InstNo <= _GEN_1599;
      end
    end else begin
      PALU0_bits_DecodeIn_InstNo <= _GEN_1599;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_DecodeIn_InstFlag <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (secondidx) begin // @[SIMDU.scala 550:32]
          PALU0_bits_DecodeIn_InstFlag <= io_DecodeIn_1_InstFlag; // @[SIMDU.scala 550:32]
        end else begin
          PALU0_bits_DecodeIn_InstFlag <= io_DecodeIn_0_InstFlag;
        end
      end else begin
        PALU0_bits_DecodeIn_InstFlag <= _GEN_1598;
      end
    end else begin
      PALU0_bits_DecodeIn_InstFlag <= _GEN_1598;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_64 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_64 <= PIDU0_io_Pctrl_isAdd_64;
        end else begin
          PALU0_bits_Pctrl_isAdd_64 <= PIDU1_io_Pctrl_isAdd_64;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_64 <= _GEN_1775;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_64 <= _GEN_1775;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_32 <= PIDU0_io_Pctrl_isAdd_32;
        end else begin
          PALU0_bits_Pctrl_isAdd_32 <= PIDU1_io_Pctrl_isAdd_32;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_32 <= _GEN_1774;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_32 <= _GEN_1774;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_16 <= PIDU0_io_Pctrl_isAdd_16;
        end else begin
          PALU0_bits_Pctrl_isAdd_16 <= PIDU1_io_Pctrl_isAdd_16;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_16 <= _GEN_1773;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_16 <= _GEN_1773;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_8 <= PIDU0_io_Pctrl_isAdd_8;
        end else begin
          PALU0_bits_Pctrl_isAdd_8 <= PIDU1_io_Pctrl_isAdd_8;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_8 <= _GEN_1772;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_8 <= _GEN_1772;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_Q15 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_Q15 <= PIDU0_io_Pctrl_isAdd_Q15;
        end else begin
          PALU0_bits_Pctrl_isAdd_Q15 <= PIDU1_io_Pctrl_isAdd_Q15;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_Q15 <= _GEN_1771;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_Q15 <= _GEN_1771;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_Q31 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_Q31 <= PIDU0_io_Pctrl_isAdd_Q31;
        end else begin
          PALU0_bits_Pctrl_isAdd_Q31 <= PIDU1_io_Pctrl_isAdd_Q31;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_Q31 <= _GEN_1770;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_Q31 <= _GEN_1770;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdd_C31 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdd_C31 <= PIDU0_io_Pctrl_isAdd_C31;
        end else begin
          PALU0_bits_Pctrl_isAdd_C31 <= PIDU1_io_Pctrl_isAdd_C31;
        end
      end else begin
        PALU0_bits_Pctrl_isAdd_C31 <= _GEN_1769;
      end
    end else begin
      PALU0_bits_Pctrl_isAdd_C31 <= _GEN_1769;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAve <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAve <= PIDU0_io_Pctrl_isAve;
        end else begin
          PALU0_bits_Pctrl_isAve <= PIDU1_io_Pctrl_isAve;
        end
      end else begin
        PALU0_bits_Pctrl_isAve <= _GEN_1768;
      end
    end else begin
      PALU0_bits_Pctrl_isAve <= _GEN_1768;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_64 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_64 <= PIDU0_io_Pctrl_isSub_64;
        end else begin
          PALU0_bits_Pctrl_isSub_64 <= PIDU1_io_Pctrl_isSub_64;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_64 <= _GEN_1766;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_64 <= _GEN_1766;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_32 <= PIDU0_io_Pctrl_isSub_32;
        end else begin
          PALU0_bits_Pctrl_isSub_32 <= PIDU1_io_Pctrl_isSub_32;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_32 <= _GEN_1765;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_32 <= _GEN_1765;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_16 <= PIDU0_io_Pctrl_isSub_16;
        end else begin
          PALU0_bits_Pctrl_isSub_16 <= PIDU1_io_Pctrl_isSub_16;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_16 <= _GEN_1764;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_16 <= _GEN_1764;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_8 <= PIDU0_io_Pctrl_isSub_8;
        end else begin
          PALU0_bits_Pctrl_isSub_8 <= PIDU1_io_Pctrl_isSub_8;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_8 <= _GEN_1763;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_8 <= _GEN_1763;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_Q15 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_Q15 <= PIDU0_io_Pctrl_isSub_Q15;
        end else begin
          PALU0_bits_Pctrl_isSub_Q15 <= PIDU1_io_Pctrl_isSub_Q15;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_Q15 <= _GEN_1762;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_Q15 <= _GEN_1762;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_Q31 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_Q31 <= PIDU0_io_Pctrl_isSub_Q31;
        end else begin
          PALU0_bits_Pctrl_isSub_Q31 <= PIDU1_io_Pctrl_isSub_Q31;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_Q31 <= _GEN_1761;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_Q31 <= _GEN_1761;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub_C31 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub_C31 <= PIDU0_io_Pctrl_isSub_C31;
        end else begin
          PALU0_bits_Pctrl_isSub_C31 <= PIDU1_io_Pctrl_isSub_C31;
        end
      end else begin
        PALU0_bits_Pctrl_isSub_C31 <= _GEN_1760;
      end
    end else begin
      PALU0_bits_Pctrl_isSub_C31 <= _GEN_1760;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCras_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCras_16 <= PIDU0_io_Pctrl_isCras_16;
        end else begin
          PALU0_bits_Pctrl_isCras_16 <= PIDU1_io_Pctrl_isCras_16;
        end
      end else begin
        PALU0_bits_Pctrl_isCras_16 <= _GEN_1759;
      end
    end else begin
      PALU0_bits_Pctrl_isCras_16 <= _GEN_1759;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCrsa_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCrsa_16 <= PIDU0_io_Pctrl_isCrsa_16;
        end else begin
          PALU0_bits_Pctrl_isCrsa_16 <= PIDU1_io_Pctrl_isCrsa_16;
        end
      end else begin
        PALU0_bits_Pctrl_isCrsa_16 <= _GEN_1758;
      end
    end else begin
      PALU0_bits_Pctrl_isCrsa_16 <= _GEN_1758;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCras_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCras_32 <= PIDU0_io_Pctrl_isCras_32;
        end else begin
          PALU0_bits_Pctrl_isCras_32 <= PIDU1_io_Pctrl_isCras_32;
        end
      end else begin
        PALU0_bits_Pctrl_isCras_32 <= _GEN_1757;
      end
    end else begin
      PALU0_bits_Pctrl_isCras_32 <= _GEN_1757;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCrsa_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCrsa_32 <= PIDU0_io_Pctrl_isCrsa_32;
        end else begin
          PALU0_bits_Pctrl_isCrsa_32 <= PIDU1_io_Pctrl_isCrsa_32;
        end
      end else begin
        PALU0_bits_Pctrl_isCrsa_32 <= _GEN_1756;
      end
    end else begin
      PALU0_bits_Pctrl_isCrsa_32 <= _GEN_1756;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isStas_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isStas_16 <= PIDU0_io_Pctrl_isStas_16;
        end else begin
          PALU0_bits_Pctrl_isStas_16 <= PIDU1_io_Pctrl_isStas_16;
        end
      end else begin
        PALU0_bits_Pctrl_isStas_16 <= _GEN_1754;
      end
    end else begin
      PALU0_bits_Pctrl_isStas_16 <= _GEN_1754;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isStsa_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isStsa_16 <= PIDU0_io_Pctrl_isStsa_16;
        end else begin
          PALU0_bits_Pctrl_isStsa_16 <= PIDU1_io_Pctrl_isStsa_16;
        end
      end else begin
        PALU0_bits_Pctrl_isStsa_16 <= _GEN_1753;
      end
    end else begin
      PALU0_bits_Pctrl_isStsa_16 <= _GEN_1753;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isStas_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isStas_32 <= PIDU0_io_Pctrl_isStas_32;
        end else begin
          PALU0_bits_Pctrl_isStas_32 <= PIDU1_io_Pctrl_isStas_32;
        end
      end else begin
        PALU0_bits_Pctrl_isStas_32 <= _GEN_1752;
      end
    end else begin
      PALU0_bits_Pctrl_isStas_32 <= _GEN_1752;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isStsa_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isStsa_32 <= PIDU0_io_Pctrl_isStsa_32;
        end else begin
          PALU0_bits_Pctrl_isStsa_32 <= PIDU1_io_Pctrl_isStsa_32;
        end
      end else begin
        PALU0_bits_Pctrl_isStsa_32 <= _GEN_1751;
      end
    end else begin
      PALU0_bits_Pctrl_isStsa_32 <= _GEN_1751;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isComp_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isComp_16 <= PIDU0_io_Pctrl_isComp_16;
        end else begin
          PALU0_bits_Pctrl_isComp_16 <= PIDU1_io_Pctrl_isComp_16;
        end
      end else begin
        PALU0_bits_Pctrl_isComp_16 <= _GEN_1749;
      end
    end else begin
      PALU0_bits_Pctrl_isComp_16 <= _GEN_1749;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isComp_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isComp_8 <= PIDU0_io_Pctrl_isComp_8;
        end else begin
          PALU0_bits_Pctrl_isComp_8 <= PIDU1_io_Pctrl_isComp_8;
        end
      end else begin
        PALU0_bits_Pctrl_isComp_8 <= _GEN_1748;
      end
    end else begin
      PALU0_bits_Pctrl_isComp_8 <= _GEN_1748;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCompare <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCompare <= PIDU0_io_Pctrl_isCompare;
        end else begin
          PALU0_bits_Pctrl_isCompare <= PIDU1_io_Pctrl_isCompare;
        end
      end else begin
        PALU0_bits_Pctrl_isCompare <= _GEN_1747;
      end
    end else begin
      PALU0_bits_Pctrl_isCompare <= _GEN_1747;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isMaxMin_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isMaxMin_16 <= PIDU0_io_Pctrl_isMaxMin_16;
        end else begin
          PALU0_bits_Pctrl_isMaxMin_16 <= PIDU1_io_Pctrl_isMaxMin_16;
        end
      end else begin
        PALU0_bits_Pctrl_isMaxMin_16 <= _GEN_1746;
      end
    end else begin
      PALU0_bits_Pctrl_isMaxMin_16 <= _GEN_1746;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isMaxMin_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isMaxMin_8 <= PIDU0_io_Pctrl_isMaxMin_8;
        end else begin
          PALU0_bits_Pctrl_isMaxMin_8 <= PIDU1_io_Pctrl_isMaxMin_8;
        end
      end else begin
        PALU0_bits_Pctrl_isMaxMin_8 <= _GEN_1745;
      end
    end else begin
      PALU0_bits_Pctrl_isMaxMin_8 <= _GEN_1745;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isMaxMin_XLEN <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isMaxMin_XLEN <= PIDU0_io_Pctrl_isMaxMin_XLEN;
        end else begin
          PALU0_bits_Pctrl_isMaxMin_XLEN <= PIDU1_io_Pctrl_isMaxMin_XLEN;
        end
      end else begin
        PALU0_bits_Pctrl_isMaxMin_XLEN <= _GEN_1744;
      end
    end else begin
      PALU0_bits_Pctrl_isMaxMin_XLEN <= _GEN_1744;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isMaxMin_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isMaxMin_32 <= PIDU0_io_Pctrl_isMaxMin_32;
        end else begin
          PALU0_bits_Pctrl_isMaxMin_32 <= PIDU1_io_Pctrl_isMaxMin_32;
        end
      end else begin
        PALU0_bits_Pctrl_isMaxMin_32 <= _GEN_1743;
      end
    end else begin
      PALU0_bits_Pctrl_isMaxMin_32 <= _GEN_1743;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isMaxMin <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isMaxMin <= PIDU0_io_Pctrl_isMaxMin;
        end else begin
          PALU0_bits_Pctrl_isMaxMin <= PIDU1_io_Pctrl_isMaxMin;
        end
      end else begin
        PALU0_bits_Pctrl_isMaxMin <= _GEN_1742;
      end
    end else begin
      PALU0_bits_Pctrl_isMaxMin <= _GEN_1742;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isPbs <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isPbs <= PIDU0_io_Pctrl_isPbs;
        end else begin
          PALU0_bits_Pctrl_isPbs <= PIDU1_io_Pctrl_isPbs;
        end
      end else begin
        PALU0_bits_Pctrl_isPbs <= _GEN_1741;
      end
    end else begin
      PALU0_bits_Pctrl_isPbs <= _GEN_1741;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isRs_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isRs_16 <= PIDU0_io_Pctrl_isRs_16;
        end else begin
          PALU0_bits_Pctrl_isRs_16 <= PIDU1_io_Pctrl_isRs_16;
        end
      end else begin
        PALU0_bits_Pctrl_isRs_16 <= _GEN_1740;
      end
    end else begin
      PALU0_bits_Pctrl_isRs_16 <= _GEN_1740;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLs_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLs_16 <= PIDU0_io_Pctrl_isLs_16;
        end else begin
          PALU0_bits_Pctrl_isLs_16 <= PIDU1_io_Pctrl_isLs_16;
        end
      end else begin
        PALU0_bits_Pctrl_isLs_16 <= _GEN_1739;
      end
    end else begin
      PALU0_bits_Pctrl_isLs_16 <= _GEN_1739;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLR_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLR_16 <= PIDU0_io_Pctrl_isLR_16;
        end else begin
          PALU0_bits_Pctrl_isLR_16 <= PIDU1_io_Pctrl_isLR_16;
        end
      end else begin
        PALU0_bits_Pctrl_isLR_16 <= _GEN_1738;
      end
    end else begin
      PALU0_bits_Pctrl_isLR_16 <= _GEN_1738;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isRs_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isRs_8 <= PIDU0_io_Pctrl_isRs_8;
        end else begin
          PALU0_bits_Pctrl_isRs_8 <= PIDU1_io_Pctrl_isRs_8;
        end
      end else begin
        PALU0_bits_Pctrl_isRs_8 <= _GEN_1737;
      end
    end else begin
      PALU0_bits_Pctrl_isRs_8 <= _GEN_1737;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLs_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLs_8 <= PIDU0_io_Pctrl_isLs_8;
        end else begin
          PALU0_bits_Pctrl_isLs_8 <= PIDU1_io_Pctrl_isLs_8;
        end
      end else begin
        PALU0_bits_Pctrl_isLs_8 <= _GEN_1736;
      end
    end else begin
      PALU0_bits_Pctrl_isLs_8 <= _GEN_1736;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLR_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLR_8 <= PIDU0_io_Pctrl_isLR_8;
        end else begin
          PALU0_bits_Pctrl_isLR_8 <= PIDU1_io_Pctrl_isLR_8;
        end
      end else begin
        PALU0_bits_Pctrl_isLR_8 <= _GEN_1735;
      end
    end else begin
      PALU0_bits_Pctrl_isLR_8 <= _GEN_1735;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isRs_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isRs_32 <= PIDU0_io_Pctrl_isRs_32;
        end else begin
          PALU0_bits_Pctrl_isRs_32 <= PIDU1_io_Pctrl_isRs_32;
        end
      end else begin
        PALU0_bits_Pctrl_isRs_32 <= _GEN_1734;
      end
    end else begin
      PALU0_bits_Pctrl_isRs_32 <= _GEN_1734;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLs_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLs_32 <= PIDU0_io_Pctrl_isLs_32;
        end else begin
          PALU0_bits_Pctrl_isLs_32 <= PIDU1_io_Pctrl_isLs_32;
        end
      end else begin
        PALU0_bits_Pctrl_isLs_32 <= _GEN_1733;
      end
    end else begin
      PALU0_bits_Pctrl_isLs_32 <= _GEN_1733;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLR_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLR_32 <= PIDU0_io_Pctrl_isLR_32;
        end else begin
          PALU0_bits_Pctrl_isLR_32 <= PIDU1_io_Pctrl_isLR_32;
        end
      end else begin
        PALU0_bits_Pctrl_isLR_32 <= _GEN_1732;
      end
    end else begin
      PALU0_bits_Pctrl_isLR_32 <= _GEN_1732;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLR_Q31 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLR_Q31 <= PIDU0_io_Pctrl_isLR_Q31;
        end else begin
          PALU0_bits_Pctrl_isLR_Q31 <= PIDU1_io_Pctrl_isLR_Q31;
        end
      end else begin
        PALU0_bits_Pctrl_isLR_Q31 <= _GEN_1731;
      end
    end else begin
      PALU0_bits_Pctrl_isLR_Q31 <= _GEN_1731;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isLs_Q31 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isLs_Q31 <= PIDU0_io_Pctrl_isLs_Q31;
        end else begin
          PALU0_bits_Pctrl_isLs_Q31 <= PIDU1_io_Pctrl_isLs_Q31;
        end
      end else begin
        PALU0_bits_Pctrl_isLs_Q31 <= _GEN_1730;
      end
    end else begin
      PALU0_bits_Pctrl_isLs_Q31 <= _GEN_1730;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isRs_XLEN <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isRs_XLEN <= PIDU0_io_Pctrl_isRs_XLEN;
        end else begin
          PALU0_bits_Pctrl_isRs_XLEN <= PIDU1_io_Pctrl_isRs_XLEN;
        end
      end else begin
        PALU0_bits_Pctrl_isRs_XLEN <= _GEN_1729;
      end
    end else begin
      PALU0_bits_Pctrl_isRs_XLEN <= _GEN_1729;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSRAIWU <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSRAIWU <= PIDU0_io_Pctrl_isSRAIWU;
        end else begin
          PALU0_bits_Pctrl_isSRAIWU <= PIDU1_io_Pctrl_isSRAIWU;
        end
      end else begin
        PALU0_bits_Pctrl_isSRAIWU <= _GEN_1728;
      end
    end else begin
      PALU0_bits_Pctrl_isSRAIWU <= _GEN_1728;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isFSRW <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isFSRW <= PIDU0_io_Pctrl_isFSRW;
        end else begin
          PALU0_bits_Pctrl_isFSRW <= PIDU1_io_Pctrl_isFSRW;
        end
      end else begin
        PALU0_bits_Pctrl_isFSRW <= _GEN_1727;
      end
    end else begin
      PALU0_bits_Pctrl_isFSRW <= _GEN_1727;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isWext <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isWext <= PIDU0_io_Pctrl_isWext;
        end else begin
          PALU0_bits_Pctrl_isWext <= PIDU1_io_Pctrl_isWext;
        end
      end else begin
        PALU0_bits_Pctrl_isWext <= _GEN_1726;
      end
    end else begin
      PALU0_bits_Pctrl_isWext <= _GEN_1726;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isShifter <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isShifter <= PIDU0_io_Pctrl_isShifter;
        end else begin
          PALU0_bits_Pctrl_isShifter <= PIDU1_io_Pctrl_isShifter;
        end
      end else begin
        PALU0_bits_Pctrl_isShifter <= _GEN_1725;
      end
    end else begin
      PALU0_bits_Pctrl_isShifter <= _GEN_1725;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isClip_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isClip_16 <= PIDU0_io_Pctrl_isClip_16;
        end else begin
          PALU0_bits_Pctrl_isClip_16 <= PIDU1_io_Pctrl_isClip_16;
        end
      end else begin
        PALU0_bits_Pctrl_isClip_16 <= _GEN_1724;
      end
    end else begin
      PALU0_bits_Pctrl_isClip_16 <= _GEN_1724;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isClip_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isClip_8 <= PIDU0_io_Pctrl_isClip_8;
        end else begin
          PALU0_bits_Pctrl_isClip_8 <= PIDU1_io_Pctrl_isClip_8;
        end
      end else begin
        PALU0_bits_Pctrl_isClip_8 <= _GEN_1723;
      end
    end else begin
      PALU0_bits_Pctrl_isClip_8 <= _GEN_1723;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isclip_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isclip_32 <= PIDU0_io_Pctrl_isclip_32;
        end else begin
          PALU0_bits_Pctrl_isclip_32 <= PIDU1_io_Pctrl_isclip_32;
        end
      end else begin
        PALU0_bits_Pctrl_isclip_32 <= _GEN_1722;
      end
    end else begin
      PALU0_bits_Pctrl_isclip_32 <= _GEN_1722;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isClip <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isClip <= PIDU0_io_Pctrl_isClip;
        end else begin
          PALU0_bits_Pctrl_isClip <= PIDU1_io_Pctrl_isClip;
        end
      end else begin
        PALU0_bits_Pctrl_isClip <= _GEN_1721;
      end
    end else begin
      PALU0_bits_Pctrl_isClip <= _GEN_1721;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSat_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSat_16 <= PIDU0_io_Pctrl_isSat_16;
        end else begin
          PALU0_bits_Pctrl_isSat_16 <= PIDU1_io_Pctrl_isSat_16;
        end
      end else begin
        PALU0_bits_Pctrl_isSat_16 <= _GEN_1720;
      end
    end else begin
      PALU0_bits_Pctrl_isSat_16 <= _GEN_1720;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSat_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSat_8 <= PIDU0_io_Pctrl_isSat_8;
        end else begin
          PALU0_bits_Pctrl_isSat_8 <= PIDU1_io_Pctrl_isSat_8;
        end
      end else begin
        PALU0_bits_Pctrl_isSat_8 <= _GEN_1719;
      end
    end else begin
      PALU0_bits_Pctrl_isSat_8 <= _GEN_1719;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSat_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSat_32 <= PIDU0_io_Pctrl_isSat_32;
        end else begin
          PALU0_bits_Pctrl_isSat_32 <= PIDU1_io_Pctrl_isSat_32;
        end
      end else begin
        PALU0_bits_Pctrl_isSat_32 <= _GEN_1718;
      end
    end else begin
      PALU0_bits_Pctrl_isSat_32 <= _GEN_1718;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSat_W <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSat_W <= PIDU0_io_Pctrl_isSat_W;
        end else begin
          PALU0_bits_Pctrl_isSat_W <= PIDU1_io_Pctrl_isSat_W;
        end
      end else begin
        PALU0_bits_Pctrl_isSat_W <= _GEN_1717;
      end
    end else begin
      PALU0_bits_Pctrl_isSat_W <= _GEN_1717;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSat <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSat <= PIDU0_io_Pctrl_isSat;
        end else begin
          PALU0_bits_Pctrl_isSat <= PIDU1_io_Pctrl_isSat;
        end
      end else begin
        PALU0_bits_Pctrl_isSat <= _GEN_1716;
      end
    end else begin
      PALU0_bits_Pctrl_isSat <= _GEN_1716;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCnt_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCnt_16 <= PIDU0_io_Pctrl_isCnt_16;
        end else begin
          PALU0_bits_Pctrl_isCnt_16 <= PIDU1_io_Pctrl_isCnt_16;
        end
      end else begin
        PALU0_bits_Pctrl_isCnt_16 <= _GEN_1715;
      end
    end else begin
      PALU0_bits_Pctrl_isCnt_16 <= _GEN_1715;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCnt_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCnt_8 <= PIDU0_io_Pctrl_isCnt_8;
        end else begin
          PALU0_bits_Pctrl_isCnt_8 <= PIDU1_io_Pctrl_isCnt_8;
        end
      end else begin
        PALU0_bits_Pctrl_isCnt_8 <= _GEN_1714;
      end
    end else begin
      PALU0_bits_Pctrl_isCnt_8 <= _GEN_1714;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCnt_32 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCnt_32 <= PIDU0_io_Pctrl_isCnt_32;
        end else begin
          PALU0_bits_Pctrl_isCnt_32 <= PIDU1_io_Pctrl_isCnt_32;
        end
      end else begin
        PALU0_bits_Pctrl_isCnt_32 <= _GEN_1713;
      end
    end else begin
      PALU0_bits_Pctrl_isCnt_32 <= _GEN_1713;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCnt <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCnt <= PIDU0_io_Pctrl_isCnt;
        end else begin
          PALU0_bits_Pctrl_isCnt <= PIDU1_io_Pctrl_isCnt;
        end
      end else begin
        PALU0_bits_Pctrl_isCnt <= _GEN_1712;
      end
    end else begin
      PALU0_bits_Pctrl_isCnt <= _GEN_1712;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSwap_16 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSwap_16 <= PIDU0_io_Pctrl_isSwap_16;
        end else begin
          PALU0_bits_Pctrl_isSwap_16 <= PIDU1_io_Pctrl_isSwap_16;
        end
      end else begin
        PALU0_bits_Pctrl_isSwap_16 <= _GEN_1711;
      end
    end else begin
      PALU0_bits_Pctrl_isSwap_16 <= _GEN_1711;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSwap_8 <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSwap_8 <= PIDU0_io_Pctrl_isSwap_8;
        end else begin
          PALU0_bits_Pctrl_isSwap_8 <= PIDU1_io_Pctrl_isSwap_8;
        end
      end else begin
        PALU0_bits_Pctrl_isSwap_8 <= _GEN_1710;
      end
    end else begin
      PALU0_bits_Pctrl_isSwap_8 <= _GEN_1710;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSwap <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSwap <= PIDU0_io_Pctrl_isSwap;
        end else begin
          PALU0_bits_Pctrl_isSwap <= PIDU1_io_Pctrl_isSwap;
        end
      end else begin
        PALU0_bits_Pctrl_isSwap <= _GEN_1709;
      end
    end else begin
      PALU0_bits_Pctrl_isSwap <= _GEN_1709;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isUnpack <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isUnpack <= PIDU0_io_Pctrl_isUnpack;
        end else begin
          PALU0_bits_Pctrl_isUnpack <= PIDU1_io_Pctrl_isUnpack;
        end
      end else begin
        PALU0_bits_Pctrl_isUnpack <= _GEN_1708;
      end
    end else begin
      PALU0_bits_Pctrl_isUnpack <= _GEN_1708;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isBitrev <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isBitrev <= PIDU0_io_Pctrl_isBitrev;
        end else begin
          PALU0_bits_Pctrl_isBitrev <= PIDU1_io_Pctrl_isBitrev;
        end
      end else begin
        PALU0_bits_Pctrl_isBitrev <= _GEN_1707;
      end
    end else begin
      PALU0_bits_Pctrl_isBitrev <= _GEN_1707;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isCmix <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isCmix <= PIDU0_io_Pctrl_isCmix;
        end else begin
          PALU0_bits_Pctrl_isCmix <= PIDU1_io_Pctrl_isCmix;
        end
      end else begin
        PALU0_bits_Pctrl_isCmix <= _GEN_1706;
      end
    end else begin
      PALU0_bits_Pctrl_isCmix <= _GEN_1706;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isInsertb <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isInsertb <= PIDU0_io_Pctrl_isInsertb;
        end else begin
          PALU0_bits_Pctrl_isInsertb <= PIDU1_io_Pctrl_isInsertb;
        end
      end else begin
        PALU0_bits_Pctrl_isInsertb <= _GEN_1705;
      end
    end else begin
      PALU0_bits_Pctrl_isInsertb <= _GEN_1705;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isPackbb <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isPackbb <= PIDU0_io_Pctrl_isPackbb;
        end else begin
          PALU0_bits_Pctrl_isPackbb <= PIDU1_io_Pctrl_isPackbb;
        end
      end else begin
        PALU0_bits_Pctrl_isPackbb <= _GEN_1704;
      end
    end else begin
      PALU0_bits_Pctrl_isPackbb <= _GEN_1704;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isPackbt <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isPackbt <= PIDU0_io_Pctrl_isPackbt;
        end else begin
          PALU0_bits_Pctrl_isPackbt <= PIDU1_io_Pctrl_isPackbt;
        end
      end else begin
        PALU0_bits_Pctrl_isPackbt <= _GEN_1703;
      end
    end else begin
      PALU0_bits_Pctrl_isPackbt <= _GEN_1703;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isPacktb <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isPacktb <= PIDU0_io_Pctrl_isPacktb;
        end else begin
          PALU0_bits_Pctrl_isPacktb <= PIDU1_io_Pctrl_isPacktb;
        end
      end else begin
        PALU0_bits_Pctrl_isPacktb <= _GEN_1702;
      end
    end else begin
      PALU0_bits_Pctrl_isPacktb <= _GEN_1702;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isPacktt <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isPacktt <= PIDU0_io_Pctrl_isPacktt;
        end else begin
          PALU0_bits_Pctrl_isPacktt <= PIDU1_io_Pctrl_isPacktt;
        end
      end else begin
        PALU0_bits_Pctrl_isPacktt <= _GEN_1701;
      end
    end else begin
      PALU0_bits_Pctrl_isPacktt <= _GEN_1701;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isPack <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isPack <= PIDU0_io_Pctrl_isPack;
        end else begin
          PALU0_bits_Pctrl_isPack <= PIDU1_io_Pctrl_isPack;
        end
      end else begin
        PALU0_bits_Pctrl_isPack <= _GEN_1700;
      end
    end else begin
      PALU0_bits_Pctrl_isPack <= _GEN_1700;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isSub <= 8'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isSub <= PIDU0_io_Pctrl_isSub;
        end else begin
          PALU0_bits_Pctrl_isSub <= PIDU1_io_Pctrl_isSub;
        end
      end else begin
        PALU0_bits_Pctrl_isSub <= _GEN_1699;
      end
    end else begin
      PALU0_bits_Pctrl_isSub <= _GEN_1699;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_isAdder <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_isAdder <= PIDU0_io_Pctrl_isAdder;
        end else begin
          PALU0_bits_Pctrl_isAdder <= PIDU1_io_Pctrl_isAdder;
        end
      end else begin
        PALU0_bits_Pctrl_isAdder <= _GEN_1698;
      end
    end else begin
      PALU0_bits_Pctrl_isAdder <= _GEN_1698;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_SrcSigned <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_SrcSigned <= PIDU0_io_Pctrl_SrcSigned;
        end else begin
          PALU0_bits_Pctrl_SrcSigned <= PIDU1_io_Pctrl_SrcSigned;
        end
      end else begin
        PALU0_bits_Pctrl_SrcSigned <= _GEN_1697;
      end
    end else begin
      PALU0_bits_Pctrl_SrcSigned <= _GEN_1697;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_Saturating <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_Saturating <= PIDU0_io_Pctrl_Saturating;
        end else begin
          PALU0_bits_Pctrl_Saturating <= PIDU1_io_Pctrl_Saturating;
        end
      end else begin
        PALU0_bits_Pctrl_Saturating <= _GEN_1696;
      end
    end else begin
      PALU0_bits_Pctrl_Saturating <= _GEN_1696;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_Translation <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_Translation <= PIDU0_io_Pctrl_Translation;
        end else begin
          PALU0_bits_Pctrl_Translation <= PIDU1_io_Pctrl_Translation;
        end
      end else begin
        PALU0_bits_Pctrl_Translation <= _GEN_1695;
      end
    end else begin
      PALU0_bits_Pctrl_Translation <= _GEN_1695;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_LessEqual <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_LessEqual <= PIDU0_io_Pctrl_LessEqual;
        end else begin
          PALU0_bits_Pctrl_LessEqual <= PIDU1_io_Pctrl_LessEqual;
        end
      end else begin
        PALU0_bits_Pctrl_LessEqual <= _GEN_1694;
      end
    end else begin
      PALU0_bits_Pctrl_LessEqual <= _GEN_1694;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_LessThan <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_LessThan <= PIDU0_io_Pctrl_LessThan;
        end else begin
          PALU0_bits_Pctrl_LessThan <= PIDU1_io_Pctrl_LessThan;
        end
      end else begin
        PALU0_bits_Pctrl_LessThan <= _GEN_1693;
      end
    end else begin
      PALU0_bits_Pctrl_LessThan <= _GEN_1693;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_adderRes_ori <= 80'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_adderRes_ori <= PIDU0_io_Pctrl_adderRes_ori;
        end else begin
          PALU0_bits_Pctrl_adderRes_ori <= PIDU1_io_Pctrl_adderRes_ori;
        end
      end else begin
        PALU0_bits_Pctrl_adderRes_ori <= _GEN_1692;
      end
    end else begin
      PALU0_bits_Pctrl_adderRes_ori <= _GEN_1692;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_adderRes <= 64'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_adderRes <= PIDU0_io_Pctrl_adderRes;
        end else begin
          PALU0_bits_Pctrl_adderRes <= PIDU1_io_Pctrl_adderRes;
        end
      end else begin
        PALU0_bits_Pctrl_adderRes <= _GEN_1691;
      end
    end else begin
      PALU0_bits_Pctrl_adderRes <= _GEN_1691;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_adderRes_ori_drophighestbit <= 80'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_adderRes_ori_drophighestbit <= PIDU0_io_Pctrl_adderRes_ori_drophighestbit;
        end else begin
          PALU0_bits_Pctrl_adderRes_ori_drophighestbit <= PIDU1_io_Pctrl_adderRes_ori_drophighestbit;
        end
      end else begin
        PALU0_bits_Pctrl_adderRes_ori_drophighestbit <= _GEN_1690;
      end
    end else begin
      PALU0_bits_Pctrl_adderRes_ori_drophighestbit <= _GEN_1690;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_Round <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_Round <= PIDU0_io_Pctrl_Round;
        end else begin
          PALU0_bits_Pctrl_Round <= PIDU1_io_Pctrl_Round;
        end
      end else begin
        PALU0_bits_Pctrl_Round <= _GEN_1689;
      end
    end else begin
      PALU0_bits_Pctrl_Round <= _GEN_1689;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_ShiftSigned <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_ShiftSigned <= PIDU0_io_Pctrl_ShiftSigned;
        end else begin
          PALU0_bits_Pctrl_ShiftSigned <= PIDU1_io_Pctrl_ShiftSigned;
        end
      end else begin
        PALU0_bits_Pctrl_ShiftSigned <= _GEN_1688;
      end
    end else begin
      PALU0_bits_Pctrl_ShiftSigned <= _GEN_1688;
    end
    if (reset) begin // @[SIMDU.scala 482:32]
      PALU0_bits_Pctrl_Arithmetic <= 1'h0; // @[SIMDU.scala 482:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        if (~secondidx) begin // @[SIMDU.scala 551:38]
          PALU0_bits_Pctrl_Arithmetic <= PIDU0_io_Pctrl_Arithmetic;
        end else begin
          PALU0_bits_Pctrl_Arithmetic <= PIDU1_io_Pctrl_Arithmetic;
        end
      end else begin
        PALU0_bits_Pctrl_Arithmetic <= _GEN_1687;
      end
    end else begin
      PALU0_bits_Pctrl_Arithmetic <= _GEN_1687;
    end
    if (reset) begin // @[SIMDU.scala 484:28]
      PALU0_valid <= 1'h0; // @[SIMDU.scala 484:28]
    end else if (io_flush) begin // @[SIMDU.scala 572:17]
      PALU0_valid <= 1'h0; // @[SIMDU.scala 572:35]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PALU0_valid <= _GEN_2637;
    end else if (_GEN_7 & (_GEN_5 == 5'h14 | _GEN_5 == 5'h17 | _GEN_5 == 5'h15)) begin // @[SIMDU.scala 518:180]
      PALU0_valid <= _GEN_325;
    end else begin
      PALU0_valid <= _GEN_0;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_cf_pc <= 39'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_cf_pc <= _GEN_1844;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_cf_pc <= _GEN_2449; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_cf_pc <= _GEN_1844;
      end
    end else begin
      PALU1_bits_DecodeIn_cf_pc <= _GEN_1844;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_cf_runahead_checkpoint_id <= 64'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1808;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_2377; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1808;
      end
    end else begin
      PALU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1808;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_ctrl_fuOpType <= 7'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_1802;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_2367; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_1802;
      end
    end else begin
      PALU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_1802;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_ctrl_funct3 <= 3'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_ctrl_funct3 <= _GEN_1801;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_ctrl_funct3 <= _GEN_2365; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_ctrl_funct3 <= _GEN_1801;
      end
    end else begin
      PALU1_bits_DecodeIn_ctrl_funct3 <= _GEN_1801;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_ctrl_func24 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_ctrl_func24 <= _GEN_1800;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_ctrl_func24 <= _GEN_2363; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_ctrl_func24 <= _GEN_1800;
      end
    end else begin
      PALU1_bits_DecodeIn_ctrl_func24 <= _GEN_1800;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_ctrl_rfWen <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_ctrl_rfWen <= _GEN_1795;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_ctrl_rfWen <= _GEN_2353; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_ctrl_rfWen <= _GEN_1795;
      end
    end else begin
      PALU1_bits_DecodeIn_ctrl_rfWen <= _GEN_1795;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_ctrl_rfDest <= 5'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_ctrl_rfDest <= _GEN_1794;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_ctrl_rfDest <= _GEN_2351; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_ctrl_rfDest <= _GEN_1794;
      end
    end else begin
      PALU1_bits_DecodeIn_ctrl_rfDest <= _GEN_1794;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_data_src1 <= 64'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_data_src1 <= _GEN_1786;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_data_src1 <= _GEN_2335; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_data_src1 <= _GEN_1786;
      end
    end else begin
      PALU1_bits_DecodeIn_data_src1 <= _GEN_1786;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_data_src2 <= 64'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_data_src2 <= _GEN_1785;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_data_src2 <= _GEN_2333; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_data_src2 <= _GEN_1785;
      end
    end else begin
      PALU1_bits_DecodeIn_data_src2 <= _GEN_1785;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_data_src3 <= 64'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_data_src3 <= _GEN_1784;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_data_src3 <= _GEN_2331; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_data_src3 <= _GEN_1784;
      end
    end else begin
      PALU1_bits_DecodeIn_data_src3 <= _GEN_1784;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_InstNo <= 5'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_InstNo <= _GEN_1781;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_InstNo <= _GEN_2325; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_InstNo <= _GEN_1781;
      end
    end else begin
      PALU1_bits_DecodeIn_InstNo <= _GEN_1781;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_DecodeIn_InstFlag <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_DecodeIn_InstFlag <= _GEN_1780;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_DecodeIn_InstFlag <= _GEN_2323; // @[SIMDU.scala 555:32]
      end else begin
        PALU1_bits_DecodeIn_InstFlag <= _GEN_1780;
      end
    end else begin
      PALU1_bits_DecodeIn_InstFlag <= _GEN_1780;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_64 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_64 <= _GEN_1957;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_64 <= _T_43_isAdd_64; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_64 <= _GEN_1957;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_64 <= _GEN_1957;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_32 <= _GEN_1956;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_32 <= _T_43_isAdd_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_32 <= _GEN_1956;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_32 <= _GEN_1956;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_16 <= _GEN_1955;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_16 <= _T_43_isAdd_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_16 <= _GEN_1955;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_16 <= _GEN_1955;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_8 <= _GEN_1954;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_8 <= _T_43_isAdd_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_8 <= _GEN_1954;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_8 <= _GEN_1954;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_Q15 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_Q15 <= _GEN_1953;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_Q15 <= _T_43_isAdd_Q15; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_Q15 <= _GEN_1953;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_Q15 <= _GEN_1953;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_Q31 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_Q31 <= _GEN_1952;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_Q31 <= _T_43_isAdd_Q31; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_Q31 <= _GEN_1952;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_Q31 <= _GEN_1952;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdd_C31 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdd_C31 <= _GEN_1951;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdd_C31 <= _T_43_isAdd_C31; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdd_C31 <= _GEN_1951;
      end
    end else begin
      PALU1_bits_Pctrl_isAdd_C31 <= _GEN_1951;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAve <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAve <= _GEN_1950;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAve <= _T_43_isAve; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAve <= _GEN_1950;
      end
    end else begin
      PALU1_bits_Pctrl_isAve <= _GEN_1950;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_64 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_64 <= _GEN_1948;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_64 <= _T_43_isSub_64; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_64 <= _GEN_1948;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_64 <= _GEN_1948;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_32 <= _GEN_1947;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_32 <= _T_43_isSub_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_32 <= _GEN_1947;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_32 <= _GEN_1947;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_16 <= _GEN_1946;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_16 <= _T_43_isSub_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_16 <= _GEN_1946;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_16 <= _GEN_1946;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_8 <= _GEN_1945;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_8 <= _T_43_isSub_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_8 <= _GEN_1945;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_8 <= _GEN_1945;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_Q15 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_Q15 <= _GEN_1944;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_Q15 <= _T_43_isSub_Q15; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_Q15 <= _GEN_1944;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_Q15 <= _GEN_1944;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_Q31 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_Q31 <= _GEN_1943;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_Q31 <= _T_43_isSub_Q31; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_Q31 <= _GEN_1943;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_Q31 <= _GEN_1943;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub_C31 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub_C31 <= _GEN_1942;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub_C31 <= _T_43_isSub_C31; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub_C31 <= _GEN_1942;
      end
    end else begin
      PALU1_bits_Pctrl_isSub_C31 <= _GEN_1942;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCras_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCras_16 <= _GEN_1941;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCras_16 <= _T_43_isCras_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCras_16 <= _GEN_1941;
      end
    end else begin
      PALU1_bits_Pctrl_isCras_16 <= _GEN_1941;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCrsa_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCrsa_16 <= _GEN_1940;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCrsa_16 <= _T_43_isCrsa_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCrsa_16 <= _GEN_1940;
      end
    end else begin
      PALU1_bits_Pctrl_isCrsa_16 <= _GEN_1940;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCras_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCras_32 <= _GEN_1939;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCras_32 <= _T_43_isCras_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCras_32 <= _GEN_1939;
      end
    end else begin
      PALU1_bits_Pctrl_isCras_32 <= _GEN_1939;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCrsa_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCrsa_32 <= _GEN_1938;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCrsa_32 <= _T_43_isCrsa_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCrsa_32 <= _GEN_1938;
      end
    end else begin
      PALU1_bits_Pctrl_isCrsa_32 <= _GEN_1938;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isStas_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isStas_16 <= _GEN_1936;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isStas_16 <= _T_43_isStas_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isStas_16 <= _GEN_1936;
      end
    end else begin
      PALU1_bits_Pctrl_isStas_16 <= _GEN_1936;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isStsa_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isStsa_16 <= _GEN_1935;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isStsa_16 <= _T_43_isStsa_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isStsa_16 <= _GEN_1935;
      end
    end else begin
      PALU1_bits_Pctrl_isStsa_16 <= _GEN_1935;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isStas_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isStas_32 <= _GEN_1934;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isStas_32 <= _T_43_isStas_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isStas_32 <= _GEN_1934;
      end
    end else begin
      PALU1_bits_Pctrl_isStas_32 <= _GEN_1934;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isStsa_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isStsa_32 <= _GEN_1933;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isStsa_32 <= _T_43_isStsa_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isStsa_32 <= _GEN_1933;
      end
    end else begin
      PALU1_bits_Pctrl_isStsa_32 <= _GEN_1933;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isComp_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isComp_16 <= _GEN_1931;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isComp_16 <= _T_43_isComp_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isComp_16 <= _GEN_1931;
      end
    end else begin
      PALU1_bits_Pctrl_isComp_16 <= _GEN_1931;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isComp_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isComp_8 <= _GEN_1930;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isComp_8 <= _T_43_isComp_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isComp_8 <= _GEN_1930;
      end
    end else begin
      PALU1_bits_Pctrl_isComp_8 <= _GEN_1930;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCompare <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCompare <= _GEN_1929;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCompare <= _T_43_isCompare; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCompare <= _GEN_1929;
      end
    end else begin
      PALU1_bits_Pctrl_isCompare <= _GEN_1929;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isMaxMin_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isMaxMin_16 <= _GEN_1928;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isMaxMin_16 <= _T_43_isMaxMin_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isMaxMin_16 <= _GEN_1928;
      end
    end else begin
      PALU1_bits_Pctrl_isMaxMin_16 <= _GEN_1928;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isMaxMin_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isMaxMin_8 <= _GEN_1927;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isMaxMin_8 <= _T_43_isMaxMin_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isMaxMin_8 <= _GEN_1927;
      end
    end else begin
      PALU1_bits_Pctrl_isMaxMin_8 <= _GEN_1927;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isMaxMin_XLEN <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isMaxMin_XLEN <= _GEN_1926;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isMaxMin_XLEN <= _T_43_isMaxMin_XLEN; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isMaxMin_XLEN <= _GEN_1926;
      end
    end else begin
      PALU1_bits_Pctrl_isMaxMin_XLEN <= _GEN_1926;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isMaxMin_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isMaxMin_32 <= _GEN_1925;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isMaxMin_32 <= _T_43_isMaxMin_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isMaxMin_32 <= _GEN_1925;
      end
    end else begin
      PALU1_bits_Pctrl_isMaxMin_32 <= _GEN_1925;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isMaxMin <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isMaxMin <= _GEN_1924;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isMaxMin <= _T_43_isMaxMin; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isMaxMin <= _GEN_1924;
      end
    end else begin
      PALU1_bits_Pctrl_isMaxMin <= _GEN_1924;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isPbs <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isPbs <= _GEN_1923;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isPbs <= _T_43_isPbs; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isPbs <= _GEN_1923;
      end
    end else begin
      PALU1_bits_Pctrl_isPbs <= _GEN_1923;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isRs_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isRs_16 <= _GEN_1922;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isRs_16 <= _T_43_isRs_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isRs_16 <= _GEN_1922;
      end
    end else begin
      PALU1_bits_Pctrl_isRs_16 <= _GEN_1922;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLs_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLs_16 <= _GEN_1921;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLs_16 <= _T_43_isLs_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLs_16 <= _GEN_1921;
      end
    end else begin
      PALU1_bits_Pctrl_isLs_16 <= _GEN_1921;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLR_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLR_16 <= _GEN_1920;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLR_16 <= _T_43_isLR_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLR_16 <= _GEN_1920;
      end
    end else begin
      PALU1_bits_Pctrl_isLR_16 <= _GEN_1920;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isRs_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isRs_8 <= _GEN_1919;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isRs_8 <= _T_43_isRs_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isRs_8 <= _GEN_1919;
      end
    end else begin
      PALU1_bits_Pctrl_isRs_8 <= _GEN_1919;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLs_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLs_8 <= _GEN_1918;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLs_8 <= _T_43_isLs_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLs_8 <= _GEN_1918;
      end
    end else begin
      PALU1_bits_Pctrl_isLs_8 <= _GEN_1918;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLR_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLR_8 <= _GEN_1917;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLR_8 <= _T_43_isLR_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLR_8 <= _GEN_1917;
      end
    end else begin
      PALU1_bits_Pctrl_isLR_8 <= _GEN_1917;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isRs_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isRs_32 <= _GEN_1916;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isRs_32 <= _T_43_isRs_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isRs_32 <= _GEN_1916;
      end
    end else begin
      PALU1_bits_Pctrl_isRs_32 <= _GEN_1916;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLs_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLs_32 <= _GEN_1915;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLs_32 <= _T_43_isLs_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLs_32 <= _GEN_1915;
      end
    end else begin
      PALU1_bits_Pctrl_isLs_32 <= _GEN_1915;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLR_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLR_32 <= _GEN_1914;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLR_32 <= _T_43_isLR_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLR_32 <= _GEN_1914;
      end
    end else begin
      PALU1_bits_Pctrl_isLR_32 <= _GEN_1914;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLR_Q31 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLR_Q31 <= _GEN_1913;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLR_Q31 <= _T_43_isLR_Q31; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLR_Q31 <= _GEN_1913;
      end
    end else begin
      PALU1_bits_Pctrl_isLR_Q31 <= _GEN_1913;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isLs_Q31 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isLs_Q31 <= _GEN_1912;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isLs_Q31 <= _T_43_isLs_Q31; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isLs_Q31 <= _GEN_1912;
      end
    end else begin
      PALU1_bits_Pctrl_isLs_Q31 <= _GEN_1912;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isRs_XLEN <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isRs_XLEN <= _GEN_1911;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isRs_XLEN <= _T_43_isRs_XLEN; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isRs_XLEN <= _GEN_1911;
      end
    end else begin
      PALU1_bits_Pctrl_isRs_XLEN <= _GEN_1911;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSRAIWU <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSRAIWU <= _GEN_1910;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSRAIWU <= _T_43_isSRAIWU; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSRAIWU <= _GEN_1910;
      end
    end else begin
      PALU1_bits_Pctrl_isSRAIWU <= _GEN_1910;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isFSRW <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isFSRW <= _GEN_1909;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isFSRW <= _T_43_isFSRW; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isFSRW <= _GEN_1909;
      end
    end else begin
      PALU1_bits_Pctrl_isFSRW <= _GEN_1909;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isWext <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isWext <= _GEN_1908;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isWext <= _T_43_isWext; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isWext <= _GEN_1908;
      end
    end else begin
      PALU1_bits_Pctrl_isWext <= _GEN_1908;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isShifter <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isShifter <= _GEN_1907;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isShifter <= _T_43_isShifter; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isShifter <= _GEN_1907;
      end
    end else begin
      PALU1_bits_Pctrl_isShifter <= _GEN_1907;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isClip_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isClip_16 <= _GEN_1906;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isClip_16 <= _T_43_isClip_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isClip_16 <= _GEN_1906;
      end
    end else begin
      PALU1_bits_Pctrl_isClip_16 <= _GEN_1906;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isClip_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isClip_8 <= _GEN_1905;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isClip_8 <= _T_43_isClip_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isClip_8 <= _GEN_1905;
      end
    end else begin
      PALU1_bits_Pctrl_isClip_8 <= _GEN_1905;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isclip_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isclip_32 <= _GEN_1904;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isclip_32 <= _T_43_isclip_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isclip_32 <= _GEN_1904;
      end
    end else begin
      PALU1_bits_Pctrl_isclip_32 <= _GEN_1904;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isClip <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isClip <= _GEN_1903;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isClip <= _T_43_isClip; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isClip <= _GEN_1903;
      end
    end else begin
      PALU1_bits_Pctrl_isClip <= _GEN_1903;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSat_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSat_16 <= _GEN_1902;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSat_16 <= _T_43_isSat_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSat_16 <= _GEN_1902;
      end
    end else begin
      PALU1_bits_Pctrl_isSat_16 <= _GEN_1902;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSat_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSat_8 <= _GEN_1901;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSat_8 <= _T_43_isSat_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSat_8 <= _GEN_1901;
      end
    end else begin
      PALU1_bits_Pctrl_isSat_8 <= _GEN_1901;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSat_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSat_32 <= _GEN_1900;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSat_32 <= _T_43_isSat_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSat_32 <= _GEN_1900;
      end
    end else begin
      PALU1_bits_Pctrl_isSat_32 <= _GEN_1900;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSat_W <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSat_W <= _GEN_1899;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSat_W <= _T_43_isSat_W; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSat_W <= _GEN_1899;
      end
    end else begin
      PALU1_bits_Pctrl_isSat_W <= _GEN_1899;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSat <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSat <= _GEN_1898;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSat <= _T_43_isSat; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSat <= _GEN_1898;
      end
    end else begin
      PALU1_bits_Pctrl_isSat <= _GEN_1898;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCnt_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCnt_16 <= _GEN_1897;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCnt_16 <= _T_43_isCnt_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCnt_16 <= _GEN_1897;
      end
    end else begin
      PALU1_bits_Pctrl_isCnt_16 <= _GEN_1897;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCnt_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCnt_8 <= _GEN_1896;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCnt_8 <= _T_43_isCnt_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCnt_8 <= _GEN_1896;
      end
    end else begin
      PALU1_bits_Pctrl_isCnt_8 <= _GEN_1896;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCnt_32 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCnt_32 <= _GEN_1895;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCnt_32 <= _T_43_isCnt_32; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCnt_32 <= _GEN_1895;
      end
    end else begin
      PALU1_bits_Pctrl_isCnt_32 <= _GEN_1895;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCnt <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCnt <= _GEN_1894;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCnt <= _T_43_isCnt; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCnt <= _GEN_1894;
      end
    end else begin
      PALU1_bits_Pctrl_isCnt <= _GEN_1894;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSwap_16 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSwap_16 <= _GEN_1893;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSwap_16 <= _T_43_isSwap_16; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSwap_16 <= _GEN_1893;
      end
    end else begin
      PALU1_bits_Pctrl_isSwap_16 <= _GEN_1893;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSwap_8 <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSwap_8 <= _GEN_1892;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSwap_8 <= _T_43_isSwap_8; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSwap_8 <= _GEN_1892;
      end
    end else begin
      PALU1_bits_Pctrl_isSwap_8 <= _GEN_1892;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSwap <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSwap <= _GEN_1891;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSwap <= _T_43_isSwap; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSwap <= _GEN_1891;
      end
    end else begin
      PALU1_bits_Pctrl_isSwap <= _GEN_1891;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isUnpack <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isUnpack <= _GEN_1890;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isUnpack <= _T_43_isUnpack; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isUnpack <= _GEN_1890;
      end
    end else begin
      PALU1_bits_Pctrl_isUnpack <= _GEN_1890;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isBitrev <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isBitrev <= _GEN_1889;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isBitrev <= _T_43_isBitrev; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isBitrev <= _GEN_1889;
      end
    end else begin
      PALU1_bits_Pctrl_isBitrev <= _GEN_1889;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isCmix <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isCmix <= _GEN_1888;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isCmix <= _T_43_isCmix; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isCmix <= _GEN_1888;
      end
    end else begin
      PALU1_bits_Pctrl_isCmix <= _GEN_1888;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isInsertb <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isInsertb <= _GEN_1887;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isInsertb <= _T_43_isInsertb; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isInsertb <= _GEN_1887;
      end
    end else begin
      PALU1_bits_Pctrl_isInsertb <= _GEN_1887;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isPackbb <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isPackbb <= _GEN_1886;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isPackbb <= _T_43_isPackbb; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isPackbb <= _GEN_1886;
      end
    end else begin
      PALU1_bits_Pctrl_isPackbb <= _GEN_1886;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isPackbt <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isPackbt <= _GEN_1885;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isPackbt <= _T_43_isPackbt; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isPackbt <= _GEN_1885;
      end
    end else begin
      PALU1_bits_Pctrl_isPackbt <= _GEN_1885;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isPacktb <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isPacktb <= _GEN_1884;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isPacktb <= _T_43_isPacktb; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isPacktb <= _GEN_1884;
      end
    end else begin
      PALU1_bits_Pctrl_isPacktb <= _GEN_1884;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isPacktt <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isPacktt <= _GEN_1883;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isPacktt <= _T_43_isPacktt; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isPacktt <= _GEN_1883;
      end
    end else begin
      PALU1_bits_Pctrl_isPacktt <= _GEN_1883;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isPack <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isPack <= _GEN_1882;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isPack <= _T_43_isPack; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isPack <= _GEN_1882;
      end
    end else begin
      PALU1_bits_Pctrl_isPack <= _GEN_1882;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isSub <= 8'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isSub <= _GEN_1881;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isSub <= _T_43_isSub; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isSub <= _GEN_1881;
      end
    end else begin
      PALU1_bits_Pctrl_isSub <= _GEN_1881;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_isAdder <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_isAdder <= _GEN_1880;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_isAdder <= _T_43_isAdder; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_isAdder <= _GEN_1880;
      end
    end else begin
      PALU1_bits_Pctrl_isAdder <= _GEN_1880;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_SrcSigned <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_SrcSigned <= _GEN_1879;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_SrcSigned <= _T_43_SrcSigned; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_SrcSigned <= _GEN_1879;
      end
    end else begin
      PALU1_bits_Pctrl_SrcSigned <= _GEN_1879;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_Saturating <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_Saturating <= _GEN_1878;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_Saturating <= _T_43_Saturating; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_Saturating <= _GEN_1878;
      end
    end else begin
      PALU1_bits_Pctrl_Saturating <= _GEN_1878;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_Translation <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_Translation <= _GEN_1877;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_Translation <= _T_43_Translation; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_Translation <= _GEN_1877;
      end
    end else begin
      PALU1_bits_Pctrl_Translation <= _GEN_1877;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_LessEqual <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_LessEqual <= _GEN_1876;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_LessEqual <= _T_43_LessEqual; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_LessEqual <= _GEN_1876;
      end
    end else begin
      PALU1_bits_Pctrl_LessEqual <= _GEN_1876;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_LessThan <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_LessThan <= _GEN_1875;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_LessThan <= _T_43_LessThan; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_LessThan <= _GEN_1875;
      end
    end else begin
      PALU1_bits_Pctrl_LessThan <= _GEN_1875;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_adderRes_ori <= 80'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_adderRes_ori <= _GEN_1874;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_adderRes_ori <= _T_43_adderRes_ori; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_adderRes_ori <= _GEN_1874;
      end
    end else begin
      PALU1_bits_Pctrl_adderRes_ori <= _GEN_1874;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_adderRes <= 64'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_adderRes <= _GEN_1873;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_adderRes <= _T_43_adderRes; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_adderRes <= _GEN_1873;
      end
    end else begin
      PALU1_bits_Pctrl_adderRes <= _GEN_1873;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_adderRes_ori_drophighestbit <= 80'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_adderRes_ori_drophighestbit <= _GEN_1872;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_adderRes_ori_drophighestbit <= _T_43_adderRes_ori_drophighestbit; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_adderRes_ori_drophighestbit <= _GEN_1872;
      end
    end else begin
      PALU1_bits_Pctrl_adderRes_ori_drophighestbit <= _GEN_1872;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_Round <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_Round <= _GEN_1871;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_Round <= _T_43_Round; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_Round <= _GEN_1871;
      end
    end else begin
      PALU1_bits_Pctrl_Round <= _GEN_1871;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_ShiftSigned <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_ShiftSigned <= _GEN_1870;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_ShiftSigned <= _T_43_ShiftSigned; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_ShiftSigned <= _GEN_1870;
      end
    end else begin
      PALU1_bits_Pctrl_ShiftSigned <= _GEN_1870;
    end
    if (reset) begin // @[SIMDU.scala 490:32]
      PALU1_bits_Pctrl_Arithmetic <= 1'h0; // @[SIMDU.scala 490:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_bits_Pctrl_Arithmetic <= _GEN_1869;
      end else if (PALU1_io_in_ready & ~match_operator_1) begin // @[SIMDU.scala 553:56]
        PALU1_bits_Pctrl_Arithmetic <= _T_43_Arithmetic; // @[SIMDU.scala 556:32]
      end else begin
        PALU1_bits_Pctrl_Arithmetic <= _GEN_1869;
      end
    end else begin
      PALU1_bits_Pctrl_Arithmetic <= _GEN_1869;
    end
    if (reset) begin // @[SIMDU.scala 492:28]
      PALU1_valid <= 1'h0; // @[SIMDU.scala 492:28]
    end else if (io_flush) begin // @[SIMDU.scala 577:17]
      PALU1_valid <= 1'h0; // @[SIMDU.scala 577:35]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      if (PALU0_io_in_ready & ~match_operator_0) begin // @[SIMDU.scala 548:50]
        PALU1_valid <= _GEN_1779;
      end else begin
        PALU1_valid <= _GEN_2456;
      end
    end else begin
      PALU1_valid <= _GEN_1779;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_cf_pc <= 39'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_cf_pc <= _GEN_2024;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_cf_pc <= _GEN_2449; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_cf_pc <= _GEN_2024;
      end
    end else begin
      PMDU0_bits_DecodeIn_cf_pc <= _GEN_2024;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id <= 64'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1988;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_2377; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1988;
      end
    end else begin
      PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_1988;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_ctrl_fuOpType <= 7'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_ctrl_fuOpType <= _GEN_1982;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_ctrl_fuOpType <= _GEN_2367; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_ctrl_fuOpType <= _GEN_1982;
      end
    end else begin
      PMDU0_bits_DecodeIn_ctrl_fuOpType <= _GEN_1982;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_ctrl_rfWen <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_ctrl_rfWen <= _GEN_1975;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_ctrl_rfWen <= _GEN_2353; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_ctrl_rfWen <= _GEN_1975;
      end
    end else begin
      PMDU0_bits_DecodeIn_ctrl_rfWen <= _GEN_1975;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_ctrl_rfDest <= 5'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_ctrl_rfDest <= _GEN_1974;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_ctrl_rfDest <= _GEN_2351; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_ctrl_rfDest <= _GEN_1974;
      end
    end else begin
      PMDU0_bits_DecodeIn_ctrl_rfDest <= _GEN_1974;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_data_src1 <= 64'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_data_src1 <= _GEN_1966;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_data_src1 <= _GEN_2335; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_data_src1 <= _GEN_1966;
      end
    end else begin
      PMDU0_bits_DecodeIn_data_src1 <= _GEN_1966;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_data_src2 <= 64'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_data_src2 <= _GEN_1965;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_data_src2 <= _GEN_2333; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_data_src2 <= _GEN_1965;
      end
    end else begin
      PMDU0_bits_DecodeIn_data_src2 <= _GEN_1965;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_data_src3 <= 64'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_data_src3 <= _GEN_1964;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_data_src3 <= _GEN_2331; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_data_src3 <= _GEN_1964;
      end
    end else begin
      PMDU0_bits_DecodeIn_data_src3 <= _GEN_1964;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_InstNo <= 5'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_InstNo <= _GEN_1961;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_InstNo <= _GEN_2325; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_InstNo <= _GEN_1961;
      end
    end else begin
      PMDU0_bits_DecodeIn_InstNo <= _GEN_1961;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_DecodeIn_InstFlag <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_DecodeIn_InstFlag <= _GEN_1960;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_DecodeIn_InstFlag <= _GEN_2323; // @[SIMDU.scala 562:32]
      end else begin
        PMDU0_bits_DecodeIn_InstFlag <= _GEN_1960;
      end
    end else begin
      PMDU0_bits_DecodeIn_InstFlag <= _GEN_1960;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isMul_16 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isMul_16 <= _GEN_2048;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isMul_16 <= _T_43_isMul_16; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isMul_16 <= _GEN_2048;
      end
    end else begin
      PMDU0_bits_Pctrl_isMul_16 <= _GEN_2048;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isMul_8 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isMul_8 <= _GEN_2047;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isMul_8 <= _T_43_isMul_8; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isMul_8 <= _GEN_2047;
      end
    end else begin
      PMDU0_bits_Pctrl_isMul_8 <= _GEN_2047;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isMSW_3232 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isMSW_3232 <= _GEN_2046;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isMSW_3232 <= _T_43_isMSW_3232; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isMSW_3232 <= _GEN_2046;
      end
    end else begin
      PMDU0_bits_Pctrl_isMSW_3232 <= _GEN_2046;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isMSW_3216 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isMSW_3216 <= _GEN_2045;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isMSW_3216 <= _T_43_isMSW_3216; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isMSW_3216 <= _GEN_2045;
      end
    end else begin
      PMDU0_bits_Pctrl_isMSW_3216 <= _GEN_2045;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isS1632 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isS1632 <= _GEN_2044;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isS1632 <= _T_43_isS1632; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isS1632 <= _GEN_2044;
      end
    end else begin
      PMDU0_bits_Pctrl_isS1632 <= _GEN_2044;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isS1664 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isS1664 <= _GEN_2043;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isS1664 <= _T_43_isS1664; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isS1664 <= _GEN_2043;
      end
    end else begin
      PMDU0_bits_Pctrl_isS1664 <= _GEN_2043;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_is832 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_is832 <= _GEN_2042;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_is832 <= _T_43_is832; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_is832 <= _GEN_2042;
      end
    end else begin
      PMDU0_bits_Pctrl_is832 <= _GEN_2042;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_is3264 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_is3264 <= _GEN_2041;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_is3264 <= _T_43_is3264; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_is3264 <= _GEN_2041;
      end
    end else begin
      PMDU0_bits_Pctrl_is3264 <= _GEN_2041;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_is1664 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_is1664 <= _GEN_2040;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_is1664 <= _T_43_is1664; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_is1664 <= _GEN_2040;
      end
    end else begin
      PMDU0_bits_Pctrl_is1664 <= _GEN_2040;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isQ15orQ31 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isQ15orQ31 <= _GEN_2039;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isQ15orQ31 <= _T_43_isQ15orQ31; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isQ15orQ31 <= _GEN_2039;
      end
    end else begin
      PMDU0_bits_Pctrl_isQ15orQ31 <= _GEN_2039;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isC31 <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isC31 <= _GEN_2038;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isC31 <= _T_43_isC31; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isC31 <= _GEN_2038;
      end
    end else begin
      PMDU0_bits_Pctrl_isC31 <= _GEN_2038;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isQ15_64ONLY <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isQ15_64ONLY <= _GEN_2037;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isQ15_64ONLY <= _T_43_isQ15_64ONLY; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isQ15_64ONLY <= _GEN_2037;
      end
    end else begin
      PMDU0_bits_Pctrl_isQ15_64ONLY <= _GEN_2037;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isQ63_64ONLY <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isQ63_64ONLY <= _GEN_2036;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isQ63_64ONLY <= _T_43_isQ63_64ONLY; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isQ63_64ONLY <= _GEN_2036;
      end
    end else begin
      PMDU0_bits_Pctrl_isQ63_64ONLY <= _GEN_2036;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isMul_32_64ONLY <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isMul_32_64ONLY <= _GEN_2035;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isMul_32_64ONLY <= _T_43_isMul_32_64ONLY; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isMul_32_64ONLY <= _GEN_2035;
      end
    end else begin
      PMDU0_bits_Pctrl_isMul_32_64ONLY <= _GEN_2035;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_isPMA_64ONLY <= 1'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_isPMA_64ONLY <= _GEN_2034;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_isPMA_64ONLY <= _T_43_isPMA_64ONLY; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_isPMA_64ONLY <= _GEN_2034;
      end
    end else begin
      PMDU0_bits_Pctrl_isPMA_64ONLY <= _GEN_2034;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres9_0 <= 18'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres9_0 <= _GEN_2033;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres9_0 <= _T_43_mulres9_0; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres9_0 <= _GEN_2033;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres9_0 <= _GEN_2033;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres9_1 <= 18'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres9_1 <= _GEN_2032;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres9_1 <= _T_43_mulres9_1; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres9_1 <= _GEN_2032;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres9_1 <= _GEN_2032;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres9_2 <= 18'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres9_2 <= _GEN_2031;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres9_2 <= _T_43_mulres9_2; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres9_2 <= _GEN_2031;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres9_2 <= _GEN_2031;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres9_3 <= 18'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres9_3 <= _GEN_2030;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres9_3 <= _T_43_mulres9_3; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres9_3 <= _GEN_2030;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres9_3 <= _GEN_2030;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres17_0 <= 34'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres17_0 <= _GEN_2029;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres17_0 <= _T_43_mulres17_0; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres17_0 <= _GEN_2029;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres17_0 <= _GEN_2029;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres17_1 <= 34'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres17_1 <= _GEN_2028;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres17_1 <= _T_43_mulres17_1; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres17_1 <= _GEN_2028;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres17_1 <= _GEN_2028;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres33_0 <= 66'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres33_0 <= _GEN_2027;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres33_0 <= _T_43_mulres33_0; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres33_0 <= _GEN_2027;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres33_0 <= _GEN_2027;
    end
    if (reset) begin // @[SIMDU.scala 499:32]
      PMDU0_bits_Pctrl_mulres65_0 <= 130'h0; // @[SIMDU.scala 499:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_bits_Pctrl_mulres65_0 <= _GEN_2026;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU0_bits_Pctrl_mulres65_0 <= _T_43_mulres65_0; // @[SIMDU.scala 563:32]
      end else begin
        PMDU0_bits_Pctrl_mulres65_0 <= _GEN_2026;
      end
    end else begin
      PMDU0_bits_Pctrl_mulres65_0 <= _GEN_2026;
    end
    if (reset) begin // @[SIMDU.scala 501:28]
      PMDU0_valid <= 1'h0; // @[SIMDU.scala 501:28]
    end else if (io_flush) begin // @[SIMDU.scala 582:17]
      PMDU0_valid <= 1'h0; // @[SIMDU.scala 582:35]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU0_valid <= _GEN_1959;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      PMDU0_valid <= _GEN_3182;
    end else begin
      PMDU0_valid <= _GEN_1959;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_cf_pc <= 39'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_cf_pc <= _GEN_2204;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_cf_pc <= _GEN_2204;
      end else begin
        PMDU1_bits_DecodeIn_cf_pc <= _GEN_3066;
      end
    end else begin
      PMDU1_bits_DecodeIn_cf_pc <= _GEN_2204;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id <= 64'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_2168;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_2168;
      end else begin
        PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_3030;
      end
    end else begin
      PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id <= _GEN_2168;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_ctrl_fuOpType <= 7'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_2162;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_2162;
      end else begin
        PMDU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_3024;
      end
    end else begin
      PMDU1_bits_DecodeIn_ctrl_fuOpType <= _GEN_2162;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_ctrl_rfWen <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_ctrl_rfWen <= _GEN_2155;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_ctrl_rfWen <= _GEN_2155;
      end else begin
        PMDU1_bits_DecodeIn_ctrl_rfWen <= _GEN_3017;
      end
    end else begin
      PMDU1_bits_DecodeIn_ctrl_rfWen <= _GEN_2155;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_ctrl_rfDest <= 5'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_ctrl_rfDest <= _GEN_2154;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_ctrl_rfDest <= _GEN_2154;
      end else begin
        PMDU1_bits_DecodeIn_ctrl_rfDest <= _GEN_3016;
      end
    end else begin
      PMDU1_bits_DecodeIn_ctrl_rfDest <= _GEN_2154;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_data_src1 <= 64'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_data_src1 <= _GEN_2146;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_data_src1 <= _GEN_2146;
      end else begin
        PMDU1_bits_DecodeIn_data_src1 <= _GEN_3008;
      end
    end else begin
      PMDU1_bits_DecodeIn_data_src1 <= _GEN_2146;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_data_src2 <= 64'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_data_src2 <= _GEN_2145;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_data_src2 <= _GEN_2145;
      end else begin
        PMDU1_bits_DecodeIn_data_src2 <= _GEN_3007;
      end
    end else begin
      PMDU1_bits_DecodeIn_data_src2 <= _GEN_2145;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_data_src3 <= 64'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_data_src3 <= _GEN_2144;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_data_src3 <= _GEN_2144;
      end else begin
        PMDU1_bits_DecodeIn_data_src3 <= _GEN_3006;
      end
    end else begin
      PMDU1_bits_DecodeIn_data_src3 <= _GEN_2144;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_InstNo <= 5'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_InstNo <= _GEN_2141;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_InstNo <= _GEN_2141;
      end else begin
        PMDU1_bits_DecodeIn_InstNo <= _GEN_3003;
      end
    end else begin
      PMDU1_bits_DecodeIn_InstNo <= _GEN_2141;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_DecodeIn_InstFlag <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_DecodeIn_InstFlag <= _GEN_2140;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_DecodeIn_InstFlag <= _GEN_2140;
      end else begin
        PMDU1_bits_DecodeIn_InstFlag <= _GEN_3002;
      end
    end else begin
      PMDU1_bits_DecodeIn_InstFlag <= _GEN_2140;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isMul_16 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isMul_16 <= _GEN_2228;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isMul_16 <= _GEN_2228;
      end else begin
        PMDU1_bits_Pctrl_isMul_16 <= _GEN_3090;
      end
    end else begin
      PMDU1_bits_Pctrl_isMul_16 <= _GEN_2228;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isMul_8 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isMul_8 <= _GEN_2227;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isMul_8 <= _GEN_2227;
      end else begin
        PMDU1_bits_Pctrl_isMul_8 <= _GEN_3089;
      end
    end else begin
      PMDU1_bits_Pctrl_isMul_8 <= _GEN_2227;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isMSW_3232 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isMSW_3232 <= _GEN_2226;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isMSW_3232 <= _GEN_2226;
      end else begin
        PMDU1_bits_Pctrl_isMSW_3232 <= _GEN_3088;
      end
    end else begin
      PMDU1_bits_Pctrl_isMSW_3232 <= _GEN_2226;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isMSW_3216 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isMSW_3216 <= _GEN_2225;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isMSW_3216 <= _GEN_2225;
      end else begin
        PMDU1_bits_Pctrl_isMSW_3216 <= _GEN_3087;
      end
    end else begin
      PMDU1_bits_Pctrl_isMSW_3216 <= _GEN_2225;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isS1632 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isS1632 <= _GEN_2224;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isS1632 <= _GEN_2224;
      end else begin
        PMDU1_bits_Pctrl_isS1632 <= _GEN_3086;
      end
    end else begin
      PMDU1_bits_Pctrl_isS1632 <= _GEN_2224;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isS1664 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isS1664 <= _GEN_2223;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isS1664 <= _GEN_2223;
      end else begin
        PMDU1_bits_Pctrl_isS1664 <= _GEN_3085;
      end
    end else begin
      PMDU1_bits_Pctrl_isS1664 <= _GEN_2223;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_is832 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_is832 <= _GEN_2222;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_is832 <= _GEN_2222;
      end else begin
        PMDU1_bits_Pctrl_is832 <= _GEN_3084;
      end
    end else begin
      PMDU1_bits_Pctrl_is832 <= _GEN_2222;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_is3264 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_is3264 <= _GEN_2221;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_is3264 <= _GEN_2221;
      end else begin
        PMDU1_bits_Pctrl_is3264 <= _GEN_3083;
      end
    end else begin
      PMDU1_bits_Pctrl_is3264 <= _GEN_2221;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_is1664 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_is1664 <= _GEN_2220;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_is1664 <= _GEN_2220;
      end else begin
        PMDU1_bits_Pctrl_is1664 <= _GEN_3082;
      end
    end else begin
      PMDU1_bits_Pctrl_is1664 <= _GEN_2220;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isQ15orQ31 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isQ15orQ31 <= _GEN_2219;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isQ15orQ31 <= _GEN_2219;
      end else begin
        PMDU1_bits_Pctrl_isQ15orQ31 <= _GEN_3081;
      end
    end else begin
      PMDU1_bits_Pctrl_isQ15orQ31 <= _GEN_2219;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isC31 <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isC31 <= _GEN_2218;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isC31 <= _GEN_2218;
      end else begin
        PMDU1_bits_Pctrl_isC31 <= _GEN_3080;
      end
    end else begin
      PMDU1_bits_Pctrl_isC31 <= _GEN_2218;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isQ15_64ONLY <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isQ15_64ONLY <= _GEN_2217;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isQ15_64ONLY <= _GEN_2217;
      end else begin
        PMDU1_bits_Pctrl_isQ15_64ONLY <= _GEN_3079;
      end
    end else begin
      PMDU1_bits_Pctrl_isQ15_64ONLY <= _GEN_2217;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isQ63_64ONLY <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isQ63_64ONLY <= _GEN_2216;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isQ63_64ONLY <= _GEN_2216;
      end else begin
        PMDU1_bits_Pctrl_isQ63_64ONLY <= _GEN_3078;
      end
    end else begin
      PMDU1_bits_Pctrl_isQ63_64ONLY <= _GEN_2216;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isMul_32_64ONLY <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isMul_32_64ONLY <= _GEN_2215;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isMul_32_64ONLY <= _GEN_2215;
      end else begin
        PMDU1_bits_Pctrl_isMul_32_64ONLY <= _GEN_3077;
      end
    end else begin
      PMDU1_bits_Pctrl_isMul_32_64ONLY <= _GEN_2215;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_isPMA_64ONLY <= 1'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_isPMA_64ONLY <= _GEN_2214;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_isPMA_64ONLY <= _GEN_2214;
      end else begin
        PMDU1_bits_Pctrl_isPMA_64ONLY <= _GEN_3076;
      end
    end else begin
      PMDU1_bits_Pctrl_isPMA_64ONLY <= _GEN_2214;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres9_0 <= 18'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres9_0 <= _GEN_2213;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres9_0 <= _GEN_2213;
      end else begin
        PMDU1_bits_Pctrl_mulres9_0 <= _GEN_3075;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres9_0 <= _GEN_2213;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres9_1 <= 18'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres9_1 <= _GEN_2212;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres9_1 <= _GEN_2212;
      end else begin
        PMDU1_bits_Pctrl_mulres9_1 <= _GEN_3074;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres9_1 <= _GEN_2212;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres9_2 <= 18'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres9_2 <= _GEN_2211;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres9_2 <= _GEN_2211;
      end else begin
        PMDU1_bits_Pctrl_mulres9_2 <= _GEN_3073;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres9_2 <= _GEN_2211;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres9_3 <= 18'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres9_3 <= _GEN_2210;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres9_3 <= _GEN_2210;
      end else begin
        PMDU1_bits_Pctrl_mulres9_3 <= _GEN_3072;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres9_3 <= _GEN_2210;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres17_0 <= 34'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres17_0 <= _GEN_2209;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres17_0 <= _GEN_2209;
      end else begin
        PMDU1_bits_Pctrl_mulres17_0 <= _GEN_3071;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres17_0 <= _GEN_2209;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres17_1 <= 34'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres17_1 <= _GEN_2208;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres17_1 <= _GEN_2208;
      end else begin
        PMDU1_bits_Pctrl_mulres17_1 <= _GEN_3070;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres17_1 <= _GEN_2208;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres33_0 <= 66'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres33_0 <= _GEN_2207;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres33_0 <= _GEN_2207;
      end else begin
        PMDU1_bits_Pctrl_mulres33_0 <= _GEN_3069;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres33_0 <= _GEN_2207;
    end
    if (reset) begin // @[SIMDU.scala 507:32]
      PMDU1_bits_Pctrl_mulres65_0 <= 130'h0; // @[SIMDU.scala 507:32]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_bits_Pctrl_mulres65_0 <= _GEN_2206;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      if (PMDU0_io_in_ready & ~match_operator_2) begin // @[SIMDU.scala 560:50]
        PMDU1_bits_Pctrl_mulres65_0 <= _GEN_2206;
      end else begin
        PMDU1_bits_Pctrl_mulres65_0 <= _GEN_3068;
      end
    end else begin
      PMDU1_bits_Pctrl_mulres65_0 <= _GEN_2206;
    end
    if (reset) begin // @[SIMDU.scala 509:28]
      PMDU1_valid <= 1'h0; // @[SIMDU.scala 509:28]
    end else if (io_flush) begin // @[SIMDU.scala 588:17]
      PMDU1_valid <= 1'h0; // @[SIMDU.scala 588:35]
    end else if (_GEN_2321 & (_GEN_2319 == 5'h14 | _GEN_2319 == 5'h17 | _GEN_2319 == 5'h15)) begin // @[SIMDU.scala 547:184]
      PMDU1_valid <= _GEN_2139;
    end else if (_GEN_2321 & (_GEN_2319 == 5'h16 | _GEN_2319 == 5'h1c)) begin // @[SIMDU.scala 559:142]
      PMDU1_valid <= _GEN_3363;
    end else begin
      PMDU1_valid <= _GEN_2139;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PALU0_bits_DecodeIn_cf_pc = _RAND_0[38:0];
  _RAND_1 = {2{`RANDOM}};
  PALU0_bits_DecodeIn_cf_runahead_checkpoint_id = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_ctrl_fuOpType = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_ctrl_funct3 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_ctrl_func24 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_ctrl_rfWen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_ctrl_rfDest = _RAND_6[4:0];
  _RAND_7 = {2{`RANDOM}};
  PALU0_bits_DecodeIn_data_src1 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  PALU0_bits_DecodeIn_data_src2 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  PALU0_bits_DecodeIn_data_src3 = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_InstNo = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  PALU0_bits_DecodeIn_InstFlag = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_64 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_32 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_16 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_8 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_Q15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_Q31 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdd_C31 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAve = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_64 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_32 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_16 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_8 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_Q15 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_Q31 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub_C31 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCras_16 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCrsa_16 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCras_32 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCrsa_32 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isStas_16 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isStsa_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isStas_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isStsa_32 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isComp_16 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isComp_8 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCompare = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isMaxMin_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isMaxMin_8 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isMaxMin_XLEN = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isMaxMin_32 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isMaxMin = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isPbs = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isRs_16 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLs_16 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLR_16 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isRs_8 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLs_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLR_8 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isRs_32 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLs_32 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLR_32 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLR_Q31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isLs_Q31 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isRs_XLEN = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSRAIWU = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isFSRW = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isWext = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isShifter = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isClip_16 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isClip_8 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isclip_32 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isClip = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSat_16 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSat_8 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSat_32 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSat_W = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSat = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCnt_16 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCnt_8 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCnt_32 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCnt = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSwap_16 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSwap_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSwap = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isUnpack = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isBitrev = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isCmix = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isInsertb = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isPackbb = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isPackbt = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isPacktb = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isPacktt = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isPack = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isSub = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  PALU0_bits_Pctrl_isAdder = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  PALU0_bits_Pctrl_SrcSigned = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  PALU0_bits_Pctrl_Saturating = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  PALU0_bits_Pctrl_Translation = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  PALU0_bits_Pctrl_LessEqual = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  PALU0_bits_Pctrl_LessThan = _RAND_91[0:0];
  _RAND_92 = {3{`RANDOM}};
  PALU0_bits_Pctrl_adderRes_ori = _RAND_92[79:0];
  _RAND_93 = {2{`RANDOM}};
  PALU0_bits_Pctrl_adderRes = _RAND_93[63:0];
  _RAND_94 = {3{`RANDOM}};
  PALU0_bits_Pctrl_adderRes_ori_drophighestbit = _RAND_94[79:0];
  _RAND_95 = {1{`RANDOM}};
  PALU0_bits_Pctrl_Round = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  PALU0_bits_Pctrl_ShiftSigned = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  PALU0_bits_Pctrl_Arithmetic = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  PALU0_valid = _RAND_98[0:0];
  _RAND_99 = {2{`RANDOM}};
  PALU1_bits_DecodeIn_cf_pc = _RAND_99[38:0];
  _RAND_100 = {2{`RANDOM}};
  PALU1_bits_DecodeIn_cf_runahead_checkpoint_id = _RAND_100[63:0];
  _RAND_101 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_ctrl_fuOpType = _RAND_101[6:0];
  _RAND_102 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_ctrl_funct3 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_ctrl_func24 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_ctrl_rfWen = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_ctrl_rfDest = _RAND_105[4:0];
  _RAND_106 = {2{`RANDOM}};
  PALU1_bits_DecodeIn_data_src1 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  PALU1_bits_DecodeIn_data_src2 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  PALU1_bits_DecodeIn_data_src3 = _RAND_108[63:0];
  _RAND_109 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_InstNo = _RAND_109[4:0];
  _RAND_110 = {1{`RANDOM}};
  PALU1_bits_DecodeIn_InstFlag = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_64 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_32 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_16 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_8 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_Q15 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_Q31 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdd_C31 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAve = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_64 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_32 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_16 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_8 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_Q15 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_Q31 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub_C31 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCras_16 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCrsa_16 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCras_32 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCrsa_32 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isStas_16 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isStsa_16 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isStas_32 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isStsa_32 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isComp_16 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isComp_8 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCompare = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isMaxMin_16 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isMaxMin_8 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isMaxMin_XLEN = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isMaxMin_32 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isMaxMin = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isPbs = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isRs_16 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLs_16 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLR_16 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isRs_8 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLs_8 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLR_8 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isRs_32 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLs_32 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLR_32 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLR_Q31 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isLs_Q31 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isRs_XLEN = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSRAIWU = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isFSRW = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isWext = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isShifter = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isClip_16 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isClip_8 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isclip_32 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isClip = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSat_16 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSat_8 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSat_32 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSat_W = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSat = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCnt_16 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCnt_8 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCnt_32 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCnt = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSwap_16 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSwap_8 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSwap = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isUnpack = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isBitrev = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isCmix = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isInsertb = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isPackbb = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isPackbt = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isPacktb = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isPacktt = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isPack = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isSub = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  PALU1_bits_Pctrl_isAdder = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  PALU1_bits_Pctrl_SrcSigned = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  PALU1_bits_Pctrl_Saturating = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  PALU1_bits_Pctrl_Translation = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  PALU1_bits_Pctrl_LessEqual = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  PALU1_bits_Pctrl_LessThan = _RAND_190[0:0];
  _RAND_191 = {3{`RANDOM}};
  PALU1_bits_Pctrl_adderRes_ori = _RAND_191[79:0];
  _RAND_192 = {2{`RANDOM}};
  PALU1_bits_Pctrl_adderRes = _RAND_192[63:0];
  _RAND_193 = {3{`RANDOM}};
  PALU1_bits_Pctrl_adderRes_ori_drophighestbit = _RAND_193[79:0];
  _RAND_194 = {1{`RANDOM}};
  PALU1_bits_Pctrl_Round = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  PALU1_bits_Pctrl_ShiftSigned = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  PALU1_bits_Pctrl_Arithmetic = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  PALU1_valid = _RAND_197[0:0];
  _RAND_198 = {2{`RANDOM}};
  PMDU0_bits_DecodeIn_cf_pc = _RAND_198[38:0];
  _RAND_199 = {2{`RANDOM}};
  PMDU0_bits_DecodeIn_cf_runahead_checkpoint_id = _RAND_199[63:0];
  _RAND_200 = {1{`RANDOM}};
  PMDU0_bits_DecodeIn_ctrl_fuOpType = _RAND_200[6:0];
  _RAND_201 = {1{`RANDOM}};
  PMDU0_bits_DecodeIn_ctrl_rfWen = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  PMDU0_bits_DecodeIn_ctrl_rfDest = _RAND_202[4:0];
  _RAND_203 = {2{`RANDOM}};
  PMDU0_bits_DecodeIn_data_src1 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  PMDU0_bits_DecodeIn_data_src2 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  PMDU0_bits_DecodeIn_data_src3 = _RAND_205[63:0];
  _RAND_206 = {1{`RANDOM}};
  PMDU0_bits_DecodeIn_InstNo = _RAND_206[4:0];
  _RAND_207 = {1{`RANDOM}};
  PMDU0_bits_DecodeIn_InstFlag = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isMul_16 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isMul_8 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isMSW_3232 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isMSW_3216 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isS1632 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isS1664 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_is832 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_is3264 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_is1664 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isQ15orQ31 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isC31 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isQ15_64ONLY = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isQ63_64ONLY = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isMul_32_64ONLY = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_isPMA_64ONLY = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_mulres9_0 = _RAND_223[17:0];
  _RAND_224 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_mulres9_1 = _RAND_224[17:0];
  _RAND_225 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_mulres9_2 = _RAND_225[17:0];
  _RAND_226 = {1{`RANDOM}};
  PMDU0_bits_Pctrl_mulres9_3 = _RAND_226[17:0];
  _RAND_227 = {2{`RANDOM}};
  PMDU0_bits_Pctrl_mulres17_0 = _RAND_227[33:0];
  _RAND_228 = {2{`RANDOM}};
  PMDU0_bits_Pctrl_mulres17_1 = _RAND_228[33:0];
  _RAND_229 = {3{`RANDOM}};
  PMDU0_bits_Pctrl_mulres33_0 = _RAND_229[65:0];
  _RAND_230 = {5{`RANDOM}};
  PMDU0_bits_Pctrl_mulres65_0 = _RAND_230[129:0];
  _RAND_231 = {1{`RANDOM}};
  PMDU0_valid = _RAND_231[0:0];
  _RAND_232 = {2{`RANDOM}};
  PMDU1_bits_DecodeIn_cf_pc = _RAND_232[38:0];
  _RAND_233 = {2{`RANDOM}};
  PMDU1_bits_DecodeIn_cf_runahead_checkpoint_id = _RAND_233[63:0];
  _RAND_234 = {1{`RANDOM}};
  PMDU1_bits_DecodeIn_ctrl_fuOpType = _RAND_234[6:0];
  _RAND_235 = {1{`RANDOM}};
  PMDU1_bits_DecodeIn_ctrl_rfWen = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  PMDU1_bits_DecodeIn_ctrl_rfDest = _RAND_236[4:0];
  _RAND_237 = {2{`RANDOM}};
  PMDU1_bits_DecodeIn_data_src1 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  PMDU1_bits_DecodeIn_data_src2 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  PMDU1_bits_DecodeIn_data_src3 = _RAND_239[63:0];
  _RAND_240 = {1{`RANDOM}};
  PMDU1_bits_DecodeIn_InstNo = _RAND_240[4:0];
  _RAND_241 = {1{`RANDOM}};
  PMDU1_bits_DecodeIn_InstFlag = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isMul_16 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isMul_8 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isMSW_3232 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isMSW_3216 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isS1632 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isS1664 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_is832 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_is3264 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_is1664 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isQ15orQ31 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isC31 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isQ15_64ONLY = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isQ63_64ONLY = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isMul_32_64ONLY = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_isPMA_64ONLY = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_mulres9_0 = _RAND_257[17:0];
  _RAND_258 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_mulres9_1 = _RAND_258[17:0];
  _RAND_259 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_mulres9_2 = _RAND_259[17:0];
  _RAND_260 = {1{`RANDOM}};
  PMDU1_bits_Pctrl_mulres9_3 = _RAND_260[17:0];
  _RAND_261 = {2{`RANDOM}};
  PMDU1_bits_Pctrl_mulres17_0 = _RAND_261[33:0];
  _RAND_262 = {2{`RANDOM}};
  PMDU1_bits_Pctrl_mulres17_1 = _RAND_262[33:0];
  _RAND_263 = {3{`RANDOM}};
  PMDU1_bits_Pctrl_mulres33_0 = _RAND_263[65:0];
  _RAND_264 = {5{`RANDOM}};
  PMDU1_bits_Pctrl_mulres65_0 = _RAND_264[129:0];
  _RAND_265 = {1{`RANDOM}};
  PMDU1_valid = _RAND_265[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [64:0]  io_in_bits_0,
  input  [64:0]  io_in_bits_1,
  input          io_out_ready,
  output         io_out_valid,
  output [129:0] io_out_bits,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[MDU.scala 58:22]
  wire  _T_4 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_1 = state == 2'h2 & _T_5 ? 2'h0 : state; // @[MDU.scala 80:48 81:11 84:11]
  wire [1:0] _GEN_3 = io_out_valid & ~_T_5 ? 2'h2 : _GEN_1; // @[MDU.scala 77:45 78:11]
  assign io_in_ready = state == 2'h0; // @[MDU.scala 66:24]
  assign io_out_valid = io_in_valid; // @[MDU.scala 65:16]
  assign io_out_bits = $signed(io_in_bits_0) * $signed(io_in_bits_1); // @[MDU.scala 64:37]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 58:22]
      state <= 2'h0; // @[MDU.scala 58:22]
    end else if (io_flush) begin // @[MDU.scala 68:17]
      state <= 2'h0; // @[MDU.scala 69:11]
    end else if (_T_4) begin // @[MDU.scala 71:27]
      state <= 2'h1; // @[MDU.scala 72:11]
    end else if (_T_5) begin // @[MDU.scala 74:28]
      state <= 2'h0; // @[MDU.scala 75:11]
    end else begin
      state <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [63:0]  io_in_bits_0,
  input  [63:0]  io_in_bits_1,
  input          io_sign,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[MDU.scala 102:22]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  newReq = state == 3'h0 & _T_1 & ~io_flush; // @[MDU.scala 103:51]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[MDU.scala 106:18]
  reg [128:0] shiftReg; // @[MDU.scala 108:21]
  wire [64:0] hi = shiftReg[128:64]; // @[MDU.scala 109:20]
  wire [63:0] lo = shiftReg[63:0]; // @[MDU.scala 110:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[MDU.scala 97:24]
  wire [63:0] _T_6 = 64'h0 - io_in_bits_0; // @[MDU.scala 98:16]
  wire [63:0] aVal = aSign ? _T_6 : io_in_bits_0; // @[MDU.scala 98:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[MDU.scala 97:24]
  wire [63:0] _T_9 = 64'h0 - io_in_bits_1; // @[MDU.scala 98:16]
  reg  aSignReg; // @[Reg.scala 15:16]
  wire  _T_12 = (aSign ^ bSign) & ~divBy0; // @[MDU.scala 115:44]
  reg  qSignReg; // @[Reg.scala 15:16]
  reg [63:0] bReg; // @[Reg.scala 15:16]
  wire [64:0] _T_13 = {aVal,1'h0}; // @[Cat.scala 30:58]
  reg [64:0] aValx2Reg; // @[Reg.scala 15:16]
  reg [5:0] value; // @[Counter.scala 60:40]
  wire [31:0] hi_1 = bReg[63:32]; // @[CircuitMath.scala 35:17]
  wire [31:0] lo_1 = bReg[31:0]; // @[CircuitMath.scala 36:17]
  wire  useHi = |hi_1; // @[CircuitMath.scala 37:22]
  wire [15:0] hi_2 = hi_1[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_2 = hi_1[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_1 = |hi_2; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_3 = hi_2[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_3 = hi_2[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_2 = |hi_3; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_4 = hi_3[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_4 = hi_3[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_3 = |hi_4; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_18 = hi_4[2] ? 2'h2 : {{1'd0}, hi_4[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_19 = hi_4[3] ? 2'h3 : _T_18; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_23 = lo_4[2] ? 2'h2 : {{1'd0}, lo_4[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_24 = lo_4[3] ? 2'h3 : _T_23; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_25 = useHi_3 ? _T_19 : _T_24; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_26 = {useHi_3,_T_25}; // @[Cat.scala 30:58]
  wire [3:0] hi_5 = lo_3[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_5 = lo_3[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_4 = |hi_5; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_30 = hi_5[2] ? 2'h2 : {{1'd0}, hi_5[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_31 = hi_5[3] ? 2'h3 : _T_30; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_35 = lo_5[2] ? 2'h2 : {{1'd0}, lo_5[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_36 = lo_5[3] ? 2'h3 : _T_35; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_37 = useHi_4 ? _T_31 : _T_36; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_38 = {useHi_4,_T_37}; // @[Cat.scala 30:58]
  wire [2:0] _T_39 = useHi_2 ? _T_26 : _T_38; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_40 = {useHi_2,_T_39}; // @[Cat.scala 30:58]
  wire [7:0] hi_6 = lo_2[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_6 = lo_2[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_5 = |hi_6; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_7 = hi_6[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_7 = hi_6[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_6 = |hi_7; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_44 = hi_7[2] ? 2'h2 : {{1'd0}, hi_7[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_45 = hi_7[3] ? 2'h3 : _T_44; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_49 = lo_7[2] ? 2'h2 : {{1'd0}, lo_7[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_50 = lo_7[3] ? 2'h3 : _T_49; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_51 = useHi_6 ? _T_45 : _T_50; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_52 = {useHi_6,_T_51}; // @[Cat.scala 30:58]
  wire [3:0] hi_8 = lo_6[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_8 = lo_6[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_7 = |hi_8; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_56 = hi_8[2] ? 2'h2 : {{1'd0}, hi_8[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_57 = hi_8[3] ? 2'h3 : _T_56; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_61 = lo_8[2] ? 2'h2 : {{1'd0}, lo_8[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_62 = lo_8[3] ? 2'h3 : _T_61; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_63 = useHi_7 ? _T_57 : _T_62; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_64 = {useHi_7,_T_63}; // @[Cat.scala 30:58]
  wire [2:0] _T_65 = useHi_5 ? _T_52 : _T_64; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_66 = {useHi_5,_T_65}; // @[Cat.scala 30:58]
  wire [3:0] _T_67 = useHi_1 ? _T_40 : _T_66; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_68 = {useHi_1,_T_67}; // @[Cat.scala 30:58]
  wire [15:0] hi_9 = lo_1[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_9 = lo_1[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_8 = |hi_9; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_10 = hi_9[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_10 = hi_9[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_9 = |hi_10; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_11 = hi_10[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_11 = hi_10[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_10 = |hi_11; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_72 = hi_11[2] ? 2'h2 : {{1'd0}, hi_11[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_73 = hi_11[3] ? 2'h3 : _T_72; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_77 = lo_11[2] ? 2'h2 : {{1'd0}, lo_11[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_78 = lo_11[3] ? 2'h3 : _T_77; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_79 = useHi_10 ? _T_73 : _T_78; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_80 = {useHi_10,_T_79}; // @[Cat.scala 30:58]
  wire [3:0] hi_12 = lo_10[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_12 = lo_10[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_11 = |hi_12; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_84 = hi_12[2] ? 2'h2 : {{1'd0}, hi_12[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_85 = hi_12[3] ? 2'h3 : _T_84; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_89 = lo_12[2] ? 2'h2 : {{1'd0}, lo_12[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_90 = lo_12[3] ? 2'h3 : _T_89; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_91 = useHi_11 ? _T_85 : _T_90; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_92 = {useHi_11,_T_91}; // @[Cat.scala 30:58]
  wire [2:0] _T_93 = useHi_9 ? _T_80 : _T_92; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_94 = {useHi_9,_T_93}; // @[Cat.scala 30:58]
  wire [7:0] hi_13 = lo_9[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_13 = lo_9[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_12 = |hi_13; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_14 = hi_13[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_14 = hi_13[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_13 = |hi_14; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_98 = hi_14[2] ? 2'h2 : {{1'd0}, hi_14[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_99 = hi_14[3] ? 2'h3 : _T_98; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_103 = lo_14[2] ? 2'h2 : {{1'd0}, lo_14[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_104 = lo_14[3] ? 2'h3 : _T_103; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_105 = useHi_13 ? _T_99 : _T_104; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_106 = {useHi_13,_T_105}; // @[Cat.scala 30:58]
  wire [3:0] hi_15 = lo_13[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_15 = lo_13[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_14 = |hi_15; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_110 = hi_15[2] ? 2'h2 : {{1'd0}, hi_15[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_111 = hi_15[3] ? 2'h3 : _T_110; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_115 = lo_15[2] ? 2'h2 : {{1'd0}, lo_15[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_116 = lo_15[3] ? 2'h3 : _T_115; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_117 = useHi_14 ? _T_111 : _T_116; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_118 = {useHi_14,_T_117}; // @[Cat.scala 30:58]
  wire [2:0] _T_119 = useHi_12 ? _T_106 : _T_118; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_120 = {useHi_12,_T_119}; // @[Cat.scala 30:58]
  wire [3:0] _T_121 = useHi_8 ? _T_94 : _T_120; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_122 = {useHi_8,_T_121}; // @[Cat.scala 30:58]
  wire [4:0] _T_123 = useHi ? _T_68 : _T_122; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_124 = {useHi,_T_123}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_21 = {{1'd0}, _T_124}; // @[MDU.scala 132:31]
  wire [6:0] _T_125 = 7'h40 | _GEN_21; // @[MDU.scala 132:31]
  wire  hi_16 = aValx2Reg[64]; // @[CircuitMath.scala 35:17]
  wire [63:0] lo_16 = aValx2Reg[63:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_15 = |hi_16; // @[CircuitMath.scala 37:22]
  wire [31:0] hi_17 = lo_16[63:32]; // @[CircuitMath.scala 35:17]
  wire [31:0] lo_17 = lo_16[31:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_16 = |hi_17; // @[CircuitMath.scala 37:22]
  wire [15:0] hi_18 = hi_17[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_18 = hi_17[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_17 = |hi_18; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_19 = hi_18[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_19 = hi_18[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_18 = |hi_19; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_20 = hi_19[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_20 = hi_19[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_19 = |hi_20; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_129 = hi_20[2] ? 2'h2 : {{1'd0}, hi_20[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_130 = hi_20[3] ? 2'h3 : _T_129; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_134 = lo_20[2] ? 2'h2 : {{1'd0}, lo_20[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_135 = lo_20[3] ? 2'h3 : _T_134; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_136 = useHi_19 ? _T_130 : _T_135; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_137 = {useHi_19,_T_136}; // @[Cat.scala 30:58]
  wire [3:0] hi_21 = lo_19[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_21 = lo_19[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_20 = |hi_21; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_141 = hi_21[2] ? 2'h2 : {{1'd0}, hi_21[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_142 = hi_21[3] ? 2'h3 : _T_141; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_146 = lo_21[2] ? 2'h2 : {{1'd0}, lo_21[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_147 = lo_21[3] ? 2'h3 : _T_146; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_148 = useHi_20 ? _T_142 : _T_147; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_149 = {useHi_20,_T_148}; // @[Cat.scala 30:58]
  wire [2:0] _T_150 = useHi_18 ? _T_137 : _T_149; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_151 = {useHi_18,_T_150}; // @[Cat.scala 30:58]
  wire [7:0] hi_22 = lo_18[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_22 = lo_18[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_21 = |hi_22; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_23 = hi_22[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_23 = hi_22[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_22 = |hi_23; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_155 = hi_23[2] ? 2'h2 : {{1'd0}, hi_23[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_156 = hi_23[3] ? 2'h3 : _T_155; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_160 = lo_23[2] ? 2'h2 : {{1'd0}, lo_23[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_161 = lo_23[3] ? 2'h3 : _T_160; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_162 = useHi_22 ? _T_156 : _T_161; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_163 = {useHi_22,_T_162}; // @[Cat.scala 30:58]
  wire [3:0] hi_24 = lo_22[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_24 = lo_22[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_23 = |hi_24; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_167 = hi_24[2] ? 2'h2 : {{1'd0}, hi_24[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_168 = hi_24[3] ? 2'h3 : _T_167; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_172 = lo_24[2] ? 2'h2 : {{1'd0}, lo_24[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_173 = lo_24[3] ? 2'h3 : _T_172; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_174 = useHi_23 ? _T_168 : _T_173; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_175 = {useHi_23,_T_174}; // @[Cat.scala 30:58]
  wire [2:0] _T_176 = useHi_21 ? _T_163 : _T_175; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_177 = {useHi_21,_T_176}; // @[Cat.scala 30:58]
  wire [3:0] _T_178 = useHi_17 ? _T_151 : _T_177; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_179 = {useHi_17,_T_178}; // @[Cat.scala 30:58]
  wire [15:0] hi_25 = lo_17[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_25 = lo_17[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_24 = |hi_25; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_26 = hi_25[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_26 = hi_25[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_25 = |hi_26; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_27 = hi_26[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_27 = hi_26[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_26 = |hi_27; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_183 = hi_27[2] ? 2'h2 : {{1'd0}, hi_27[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_184 = hi_27[3] ? 2'h3 : _T_183; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_188 = lo_27[2] ? 2'h2 : {{1'd0}, lo_27[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_189 = lo_27[3] ? 2'h3 : _T_188; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_190 = useHi_26 ? _T_184 : _T_189; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_191 = {useHi_26,_T_190}; // @[Cat.scala 30:58]
  wire [3:0] hi_28 = lo_26[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_28 = lo_26[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_27 = |hi_28; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_195 = hi_28[2] ? 2'h2 : {{1'd0}, hi_28[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_196 = hi_28[3] ? 2'h3 : _T_195; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_200 = lo_28[2] ? 2'h2 : {{1'd0}, lo_28[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_201 = lo_28[3] ? 2'h3 : _T_200; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_202 = useHi_27 ? _T_196 : _T_201; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_203 = {useHi_27,_T_202}; // @[Cat.scala 30:58]
  wire [2:0] _T_204 = useHi_25 ? _T_191 : _T_203; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_205 = {useHi_25,_T_204}; // @[Cat.scala 30:58]
  wire [7:0] hi_29 = lo_25[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_29 = lo_25[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_28 = |hi_29; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_30 = hi_29[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_30 = hi_29[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_29 = |hi_30; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_209 = hi_30[2] ? 2'h2 : {{1'd0}, hi_30[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_210 = hi_30[3] ? 2'h3 : _T_209; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_214 = lo_30[2] ? 2'h2 : {{1'd0}, lo_30[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_215 = lo_30[3] ? 2'h3 : _T_214; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_216 = useHi_29 ? _T_210 : _T_215; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_217 = {useHi_29,_T_216}; // @[Cat.scala 30:58]
  wire [3:0] hi_31 = lo_29[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_31 = lo_29[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_30 = |hi_31; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_221 = hi_31[2] ? 2'h2 : {{1'd0}, hi_31[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_222 = hi_31[3] ? 2'h3 : _T_221; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_226 = lo_31[2] ? 2'h2 : {{1'd0}, lo_31[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_227 = lo_31[3] ? 2'h3 : _T_226; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_228 = useHi_30 ? _T_222 : _T_227; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_229 = {useHi_30,_T_228}; // @[Cat.scala 30:58]
  wire [2:0] _T_230 = useHi_28 ? _T_217 : _T_229; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_231 = {useHi_28,_T_230}; // @[Cat.scala 30:58]
  wire [3:0] _T_232 = useHi_24 ? _T_205 : _T_231; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_233 = {useHi_24,_T_232}; // @[Cat.scala 30:58]
  wire [4:0] _T_234 = useHi_16 ? _T_179 : _T_233; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_235 = {useHi_16,_T_234}; // @[Cat.scala 30:58]
  wire [5:0] _T_236 = useHi_15 ? 6'h0 : _T_235; // @[CircuitMath.scala 38:21]
  wire [6:0] _T_237 = {useHi_15,_T_236}; // @[Cat.scala 30:58]
  wire [6:0] _T_239 = _T_125 - _T_237; // @[MDU.scala 132:45]
  wire [6:0] _value_T_1 = _T_239 >= 7'h3f ? 7'h3f : _T_239; // @[MDU.scala 136:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[MDU.scala 136:21]
  wire [127:0] _GEN_0 = {{63'd0}, aValx2Reg}; // @[MDU.scala 139:27]
  wire [127:0] _T_241 = _GEN_0 << value; // @[MDU.scala 139:27]
  wire [64:0] _GEN_22 = {{1'd0}, bReg}; // @[MDU.scala 142:28]
  wire  _T_243 = hi >= _GEN_22; // @[MDU.scala 142:28]
  wire [64:0] _T_245 = hi - _GEN_22; // @[MDU.scala 143:36]
  wire [64:0] _T_246 = _T_243 ? _T_245 : hi; // @[MDU.scala 143:24]
  wire [128:0] _T_248 = {_T_246[63:0],lo,_T_243}; // @[Cat.scala 30:58]
  wire  wrap = value == 6'h3f; // @[Counter.scala 72:24]
  wire [5:0] _value_T_4 = value + 6'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_4 = wrap ? 3'h4 : state; // @[MDU.scala 102:22 145:{36,44}]
  wire  _T_251 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_5 = state == 3'h4 & _T_251 ? 3'h0 : state; // @[MDU.scala 146:53 147:11 102:22]
  wire [128:0] _GEN_6 = state == 3'h3 ? _T_248 : shiftReg; // @[MDU.scala 141:37 143:14 108:21]
  wire [5:0] _GEN_7 = state == 3'h3 ? _value_T_4 : value; // @[MDU.scala 141:37 Counter.scala 76:15 60:40]
  wire [2:0] _GEN_8 = state == 3'h3 ? _GEN_4 : _GEN_5; // @[MDU.scala 141:37]
  wire [2:0] _GEN_10 = state == 3'h2 ? 3'h3 : _GEN_8; // @[MDU.scala 138:35 140:11]
  wire [5:0] _GEN_11 = state == 3'h2 ? value : _GEN_7; // @[MDU.scala 138:35 Counter.scala 60:40]
  wire [6:0] _GEN_12 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_11}; // @[MDU.scala 124:34 136:15]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, value} : _GEN_12; // @[MDU.scala 122:23 Counter.scala 60:40]
  wire [6:0] _GEN_19 = io_flush ? {{1'd0}, value} : _GEN_16; // @[MDU.scala 120:17 Counter.scala 60:40]
  wire [63:0] r = hi[64:1]; // @[MDU.scala 150:13]
  wire [63:0] _T_254 = 64'h0 - lo; // @[MDU.scala 151:28]
  wire [63:0] resQ = qSignReg ? _T_254 : lo; // @[MDU.scala 151:17]
  wire [63:0] _T_256 = 64'h0 - r; // @[MDU.scala 152:28]
  wire [63:0] resR = aSignReg ? _T_256 : r; // @[MDU.scala 152:17]
  assign io_in_ready = state == 3'h0; // @[MDU.scala 156:25]
  assign io_out_valid = state == 3'h4; // @[MDU.scala 155:39]
  assign io_out_bits = {resR,resQ}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 102:22]
      state <= 3'h0; // @[MDU.scala 102:22]
    end else if (io_flush) begin // @[MDU.scala 120:17]
      state <= 3'h0; // @[MDU.scala 121:11]
    end else if (newReq) begin // @[MDU.scala 122:23]
      state <= 3'h1; // @[MDU.scala 123:11]
    end else if (state == 3'h1) begin // @[MDU.scala 124:34]
      state <= 3'h2; // @[MDU.scala 137:11]
    end else begin
      state <= _GEN_10;
    end
    if (!(io_flush)) begin // @[MDU.scala 120:17]
      if (!(newReq)) begin // @[MDU.scala 122:23]
        if (!(state == 3'h1)) begin // @[MDU.scala 124:34]
          if (state == 3'h2) begin // @[MDU.scala 138:35]
            shiftReg <= {{1'd0}, _T_241}; // @[MDU.scala 139:14]
          end else begin
            shiftReg <= _GEN_6;
          end
        end
      end
    end
    if (newReq) begin // @[Reg.scala 16:19]
      aSignReg <= aSign; // @[Reg.scala 16:23]
    end
    if (newReq) begin // @[Reg.scala 16:19]
      qSignReg <= _T_12; // @[Reg.scala 16:23]
    end
    if (newReq) begin // @[Reg.scala 16:19]
      if (bSign) begin // @[MDU.scala 98:12]
        bReg <= _T_9;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin // @[Reg.scala 16:19]
      aValx2Reg <= _T_13; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 6'h0; // @[Counter.scala 60:40]
    end else begin
      value <= _GEN_19[5:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[MDU.scala 179:19]
  wire  mul_reset; // @[MDU.scala 179:19]
  wire  mul_io_in_ready; // @[MDU.scala 179:19]
  wire  mul_io_in_valid; // @[MDU.scala 179:19]
  wire [64:0] mul_io_in_bits_0; // @[MDU.scala 179:19]
  wire [64:0] mul_io_in_bits_1; // @[MDU.scala 179:19]
  wire  mul_io_out_ready; // @[MDU.scala 179:19]
  wire  mul_io_out_valid; // @[MDU.scala 179:19]
  wire [129:0] mul_io_out_bits; // @[MDU.scala 179:19]
  wire  mul_io_flush; // @[MDU.scala 179:19]
  wire  div_clock; // @[MDU.scala 180:19]
  wire  div_reset; // @[MDU.scala 180:19]
  wire  div_io_in_ready; // @[MDU.scala 180:19]
  wire  div_io_in_valid; // @[MDU.scala 180:19]
  wire [63:0] div_io_in_bits_0; // @[MDU.scala 180:19]
  wire [63:0] div_io_in_bits_1; // @[MDU.scala 180:19]
  wire  div_io_sign; // @[MDU.scala 180:19]
  wire  div_io_out_ready; // @[MDU.scala 180:19]
  wire  div_io_out_valid; // @[MDU.scala 180:19]
  wire [127:0] div_io_out_bits; // @[MDU.scala 180:19]
  wire  div_io_flush; // @[MDU.scala 180:19]
  wire  isDiv = io_in_bits_func[2]; // @[MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[MDU.scala 43:25]
  wire [64:0] _T_4 = {1'h0,io_in_bits_src1}; // @[Cat.scala 30:58]
  wire [64:0] _T_6 = {io_in_bits_src1[63],io_in_bits_src1}; // @[Cat.scala 30:58]
  wire  _T_10 = 2'h0 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_11 = 2'h1 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_12 = 2'h2 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_13 = 2'h3 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [64:0] _T_14 = _T_10 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_15 = _T_11 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_16 = _T_12 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_17 = _T_13 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_18 = _T_14 | _T_15; // @[Mux.scala 27:72]
  wire [64:0] _T_19 = _T_18 | _T_16; // @[Mux.scala 27:72]
  wire [64:0] _T_22 = {1'h0,io_in_bits_src2}; // @[Cat.scala 30:58]
  wire [64:0] _T_24 = {io_in_bits_src2[63],io_in_bits_src2}; // @[Cat.scala 30:58]
  wire [64:0] _T_31 = _T_10 ? _T_22 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_32 = _T_11 ? _T_24 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_33 = _T_12 ? _T_22 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_34 = _T_13 ? _T_22 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_35 = _T_31 | _T_32; // @[Mux.scala 27:72]
  wire [64:0] _T_36 = _T_35 | _T_33; // @[Mux.scala 27:72]
  wire [31:0] _T_41 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_42 = {_T_41,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_44 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_45 = isDivSign ? _T_42 : _T_44; // @[MDU.scala 199:47]
  wire [31:0] _T_50 = io_in_bits_src2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_51 = {_T_50,io_in_bits_src2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_53 = {32'h0,io_in_bits_src2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_54 = isDivSign ? _T_51 : _T_53; // @[MDU.scala 199:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[MDU.scala 206:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[MDU.scala 207:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[MDU.scala 208:16]
  wire [31:0] _T_69 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_70 = {_T_69,res[31:0]}; // @[Cat.scala 30:58]
  wire  _T_72 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[MDU.scala 211:50]
  wire  isDivReg = _T_72 ? isDiv : REG; // @[MDU.scala 211:21]
  wire  _T_82 = mul_io_out_ready & mul_io_out_valid; // @[Decoupled.scala 40:37]
  Multiplier mul ( // @[MDU.scala 179:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits),
    .io_flush(mul_io_flush)
  );
  Divider div ( // @[MDU.scala 180:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_ready(div_io_out_ready),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits),
    .io_flush(div_io_flush)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[MDU.scala 212:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[MDU.scala 213:22]
  assign io_out_bits = isW ? _T_70 : res; // @[MDU.scala 209:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[MDU.scala 203:34]
  assign mul_io_in_bits_0 = _T_19 | _T_17; // @[Mux.scala 27:72]
  assign mul_io_in_bits_1 = _T_36 | _T_34; // @[Mux.scala 27:72]
  assign mul_io_out_ready = io_out_ready; // @[MDU.scala 185:17]
  assign mul_io_flush = io_flush; // @[MDU.scala 181:16]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[MDU.scala 204:34]
  assign div_io_in_bits_0 = isW ? _T_45 : io_in_bits_src1; // @[MDU.scala 199:38]
  assign div_io_in_bits_1 = isW ? _T_54 : io_in_bits_src2; // @[MDU.scala 199:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[MDU.scala 42:39]
  assign div_io_out_ready = io_out_ready; // @[MDU.scala 185:17]
  assign div_io_flush = io_flush; // @[MDU.scala 182:16]
  always @(posedge clock) begin
    REG <= io_in_bits_func[2]; // @[MDU.scala 41:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU_2(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input  [38:0] io_cfIn_pnpc,
  input  [3:0]  io_cfIn_brIdx,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input  [63:0] io_offset,
  output        bpuUpdateReq_0_valid,
  output [38:0] bpuUpdateReq_0_pc,
  output        bpuUpdateReq_0_isMissPredict,
  output [38:0] bpuUpdateReq_0_actualTarget,
  output        bpuUpdateReq_0_actualTaken,
  output [6:0]  bpuUpdateReq_0_fuOpType,
  output [1:0]  bpuUpdateReq_0_btbType,
  output        bpuUpdateReq_0_isRVC
);
  wire  isAdderSub = ~io_in_bits_func[6]; // @[ALU.scala 94:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_in_bits_src2 ^ _T_2; // @[ALU.scala 95:33]
  wire [64:0] _T_4 = io_in_bits_src1 + _T_3; // @[ALU.scala 95:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 95:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 95:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[ALU.scala 96:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 97:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 98:28]
  wire [63:0] _T_10 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_14 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {_T_14,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_17 = 7'h25 == io_in_bits_func ? _T_10 : io_in_bits_src1; // @[Mux.scala 80:57]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[Mux.scala 80:57]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[ALU.scala 104:18]
  wire [126:0] _GEN_4 = {{63'd0}, shsrc1}; // @[ALU.scala 106:33]
  wire [126:0] _T_23 = _GEN_4 << shamt; // @[ALU.scala 106:33]
  wire [63:0] _T_25 = {63'h0,slt}; // @[Cat.scala 30:58]
  wire [63:0] _T_26 = {63'h0,sltu}; // @[Cat.scala 30:58]
  wire [63:0] _T_27 = shsrc1 >> shamt; // @[ALU.scala 110:32]
  wire [63:0] _T_28 = io_in_bits_src1 | io_in_bits_src2; // @[ALU.scala 111:30]
  wire [63:0] _T_29 = io_in_bits_src1 & io_in_bits_src2; // @[ALU.scala 112:30]
  wire [63:0] _T_30 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[ALU.scala 113:32]
  wire [63:0] _T_32 = $signed(_T_30) >>> shamt; // @[ALU.scala 113:49]
  wire [64:0] _T_34 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _T_23[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_36 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _T_25} : _T_34; // @[Mux.scala 80:57]
  wire [64:0] _T_38 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _T_26} : _T_36; // @[Mux.scala 80:57]
  wire [64:0] _T_40 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _T_38; // @[Mux.scala 80:57]
  wire [64:0] _T_42 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _T_27} : _T_40; // @[Mux.scala 80:57]
  wire [64:0] _T_44 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _T_28} : _T_42; // @[Mux.scala 80:57]
  wire [64:0] _T_46 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _T_29} : _T_44; // @[Mux.scala 80:57]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _T_32} : _T_46; // @[Mux.scala 80:57]
  wire [31:0] _T_52 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,res[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _T_53} : res; // @[ALU.scala 116:19]
  wire  _T_55 = ~(|xorRes); // @[ALU.scala 119:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[ALU.scala 70:30]
  wire  isBru = io_in_bits_func[4]; // @[ALU.scala 69:31]
  wire  _T_58 = 2'h0 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_59 = 2'h2 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = 2'h3 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_65 = _T_58 & _T_55 | _T_59 & slt | _T_60 & sltu; // @[Mux.scala 27:72]
  wire  taken = _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 126:72]
  wire [63:0] _GEN_1 = {{25'd0}, io_cfIn_pc}; // @[ALU.scala 127:41]
  wire [63:0] _T_68 = _GEN_1 + io_offset; // @[ALU.scala 127:41]
  wire [64:0] _T_69 = isBranch ? {{1'd0}, _T_68} : adderRes; // @[ALU.scala 127:19]
  wire [38:0] target = _T_69[38:0]; // @[ALU.scala 127:63]
  wire  _T_71 = ~taken & isBranch; // @[ALU.scala 128:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[ALU.scala 128:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 129:35]
  wire  _T_88 = ~isRVC; // @[ALU.scala 131:55]
  wire [38:0] _T_101 = io_cfIn_pc + 39'h2; // @[ALU.scala 132:71]
  wire [38:0] _T_103 = io_cfIn_pc + 39'h4; // @[ALU.scala 132:89]
  wire [38:0] _T_104 = isRVC ? _T_101 : _T_103; // @[ALU.scala 132:52]
  wire [24:0] _T_111 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_112 = {_T_111,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_114 = _T_112 + 64'h4; // @[ALU.scala 140:71]
  wire [63:0] _T_120 = _T_112 + 64'h2; // @[ALU.scala 140:108]
  wire [63:0] _T_121 = _T_88 ? _T_114 : _T_120; // @[ALU.scala 140:32]
  wire [64:0] _T_122 = isBru ? {{1'd0}, _T_121} : aluRes; // @[ALU.scala 140:21]
  wire  _T_141 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[ALU.scala 144:171]
  wire  _T_142 = io_in_bits_func == 7'h5a; // @[ALU.scala 144:205]
  wire  _T_143 = io_in_bits_func == 7'h5e; // @[ALU.scala 144:230]
  wire  _T_166 = 7'h5c == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_167 = 7'h5e == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_168 = 7'h58 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_169 = 7'h5a == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [1:0] _T_177 = _T_167 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_179 = _T_169 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_2 = {{1'd0}, _T_166}; // @[Mux.scala 27:72]
  wire [1:0] _T_186 = _GEN_2 | _T_177; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_168}; // @[Mux.scala 27:72]
  wire [1:0] _T_187 = _T_186 | _GEN_3; // @[Mux.scala 27:72]
  wire  _T_196 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_197 = _T_196 & isBru; // @[ALU.scala 157:39]
  wire  _T_230 = _T_197 & ~predictWrong; // @[ALU.scala 169:40]
  wire  _T_233 = _T_197 & predictWrong; // @[ALU.scala 170:40]
  wire  _T_234 = _T_230 & isBranch; // @[ALU.scala 171:33]
  wire  _T_235 = _T_233 & isBranch; // @[ALU.scala 172:33]
  wire  _T_239 = _T_230 & _T_141; // @[ALU.scala 173:33]
  wire  _T_243 = _T_233 & _T_141; // @[ALU.scala 174:33]
  wire  _T_245 = _T_230 & _T_142; // @[ALU.scala 175:33]
  wire  _T_247 = _T_233 & _T_142; // @[ALU.scala 176:33]
  wire  _T_249 = _T_230 & _T_143; // @[ALU.scala 177:33]
  wire  _T_251 = _T_233 & _T_143; // @[ALU.scala 178:33]
  wire [1:0] _WIRE_6 = _T_187 | _T_179; // @[Mux.scala 27:72]
  wire  bpuUpdateReq_valid = _T_196 & isBru; // @[ALU.scala 157:39]
  wire [38:0] bpuUpdateReq_pc = io_cfIn_pc;
  wire  bpuUpdateReq_isMissPredict = predictWrong; // @[ALU.scala 128:25]
  wire [38:0] bpuUpdateReq_actualTarget = target; // @[ALU.scala 127:63]
  wire  bpuUpdateReq_actualTaken = taken; // @[ALU.scala 126:72]
  wire [6:0] bpuUpdateReq_fuOpType = io_in_bits_func;
  wire [1:0] bpuUpdateReq_btbType = _T_187 | _T_179; // @[Mux.scala 27:72]
  wire  bpuUpdateReq_isRVC = isRVC; // @[ALU.scala 129:35]
  assign io_out_valid = io_in_valid; // @[ALU.scala 154:16]
  assign io_out_bits = _T_122[63:0]; // @[ALU.scala 140:15]
  assign io_redirect_target = _T_71 ? _T_104 : target; // @[ALU.scala 132:28]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[ALU.scala 134:39]
  assign bpuUpdateReq_0_valid = bpuUpdateReq_valid;
  assign bpuUpdateReq_0_pc = bpuUpdateReq_pc;
  assign bpuUpdateReq_0_isMissPredict = bpuUpdateReq_isMissPredict;
  assign bpuUpdateReq_0_actualTarget = bpuUpdateReq_actualTarget;
  assign bpuUpdateReq_0_actualTaken = bpuUpdateReq_actualTaken;
  assign bpuUpdateReq_0_fuOpType = bpuUpdateReq_fuOpType;
  assign bpuUpdateReq_0_btbType = _WIRE_6;
  assign bpuUpdateReq_0_isRVC = bpuUpdateReq_isRVC;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:130 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 130:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fatal; // @[ALU.scala 130:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module pipeline_lsu_stage1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [38:0] io_in_bits_Decode_cf_pc,
  input         io_in_bits_Decode_cf_exceptionVec_1,
  input         io_in_bits_Decode_cf_exceptionVec_2,
  input         io_in_bits_Decode_cf_exceptionVec_12,
  input         io_in_bits_Decode_cf_intrVec_0,
  input         io_in_bits_Decode_cf_intrVec_1,
  input         io_in_bits_Decode_cf_intrVec_2,
  input         io_in_bits_Decode_cf_intrVec_3,
  input         io_in_bits_Decode_cf_intrVec_4,
  input         io_in_bits_Decode_cf_intrVec_5,
  input         io_in_bits_Decode_cf_intrVec_6,
  input         io_in_bits_Decode_cf_intrVec_7,
  input         io_in_bits_Decode_cf_intrVec_8,
  input         io_in_bits_Decode_cf_intrVec_9,
  input         io_in_bits_Decode_cf_intrVec_10,
  input         io_in_bits_Decode_cf_intrVec_11,
  input         io_in_bits_Decode_cf_crossPageIPFFix,
  input  [63:0] io_in_bits_Decode_cf_runahead_checkpoint_id,
  input         io_in_bits_Decode_ctrl_rfWen,
  input  [4:0]  io_in_bits_Decode_ctrl_rfDest,
  input         io_in_bits_Decode_ctrl_isMou,
  input  [4:0]  io_in_bits_Decode_InstNo,
  input         io_in_bits_Decode_InstFlag,
  input  [63:0] io_in_bits_wdata,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_isMMIO,
  output        io_out_bits_loadAddrMisaligned,
  output        io_out_bits_storeAddrMisaligned,
  output [38:0] io_out_bits_Decode_cf_pc,
  output        io_out_bits_Decode_cf_exceptionVec_1,
  output        io_out_bits_Decode_cf_exceptionVec_2,
  output        io_out_bits_Decode_cf_exceptionVec_12,
  output        io_out_bits_Decode_cf_intrVec_0,
  output        io_out_bits_Decode_cf_intrVec_1,
  output        io_out_bits_Decode_cf_intrVec_2,
  output        io_out_bits_Decode_cf_intrVec_3,
  output        io_out_bits_Decode_cf_intrVec_4,
  output        io_out_bits_Decode_cf_intrVec_5,
  output        io_out_bits_Decode_cf_intrVec_6,
  output        io_out_bits_Decode_cf_intrVec_7,
  output        io_out_bits_Decode_cf_intrVec_8,
  output        io_out_bits_Decode_cf_intrVec_9,
  output        io_out_bits_Decode_cf_intrVec_10,
  output        io_out_bits_Decode_cf_intrVec_11,
  output        io_out_bits_Decode_cf_crossPageIPFFix,
  output [63:0] io_out_bits_Decode_cf_runahead_checkpoint_id,
  output        io_out_bits_Decode_ctrl_rfWen,
  output [4:0]  io_out_bits_Decode_ctrl_rfDest,
  output        io_out_bits_Decode_ctrl_isMou,
  output [4:0]  io_out_bits_Decode_InstNo,
  output        io_out_bits_Decode_InstFlag,
  output        io_out_bits_loadPF,
  output        io_out_bits_storePF,
  output [6:0]  io_out_bits_func,
  output [63:0] io_out_bits_addr,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_flush,
  input         DTLBPF,
  input         loadPF_0,
  input         lsuMMIO_0,
  input         storePF_0,
  input         DTLBENABLE,
  input         DTLBFINISH
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [63:0] exec_addr = io_in_bits_src1 + io_in_bits_src2; // @[SIMD_PipeLSU.scala 62:26]
  reg [1:0] req_state; // @[SIMD_PipeLSU.scala 124:26]
  wire  _T_151 = io_dmem_req_ready & io_dmem_req_valid; // @[Decoupled.scala 40:37]
  wire  exec_finish = req_state == 2'h2 | _T_151; // @[SIMD_PipeLSU.scala 164:21]
  reg  mmioReg; // @[SIMD_PipeLSU.scala 76:24]
  wire  isStore = io_in_valid & io_in_bits_func[3]; // @[SIMD_PipeLSU.scala 120:28]
  wire  _T_28 = ~isStore; // @[SIMD_PipeLSU.scala 121:21]
  wire  _T_32 = _T_151 & DTLBENABLE; // @[SIMD_PipeLSU.scala 128:29]
  wire [1:0] _GEN_11 = _T_151 & DTLBENABLE ? 2'h1 : req_state; // @[SIMD_PipeLSU.scala 124:26 128:{45,57}]
  wire  _T_36 = exec_finish & io_out_ready; // @[SIMD_PipeLSU.scala 129:76]
  wire [1:0] _T_37 = exec_finish & io_out_ready ? 2'h0 : 2'h2; // @[SIMD_PipeLSU.scala 129:63]
  wire [1:0] _GEN_12 = _T_151 & ~DTLBENABLE ? _T_37 : _GEN_11; // @[SIMD_PipeLSU.scala 129:{45,57}]
  wire  _T_40 = _T_32 & DTLBFINISH; // @[SIMD_PipeLSU.scala 130:43]
  wire [1:0] _GEN_13 = _T_32 & DTLBFINISH & DTLBPF ? 2'h0 : _GEN_12; // @[SIMD_PipeLSU.scala 130:{68,79}]
  wire  _T_45 = ~DTLBPF; // @[SIMD_PipeLSU.scala 131:60]
  wire [1:0] _GEN_15 = DTLBFINISH & DTLBPF ? 2'h0 : req_state; // @[SIMD_PipeLSU.scala 124:26 134:{36,48}]
  wire [1:0] _GEN_16 = DTLBFINISH & _T_45 ? _T_37 : _GEN_15; // @[SIMD_PipeLSU.scala 135:{36,48}]
  wire [1:0] _GEN_17 = _T_36 ? 2'h0 : req_state; // @[SIMD_PipeLSU.scala 124:26 137:{55,66}]
  wire [1:0] _GEN_18 = 2'h2 == req_state ? _GEN_17 : req_state; // @[SIMD_PipeLSU.scala 126:22 124:26]
  wire [63:0] _T_89 = {io_in_bits_wdata[7:0],io_in_bits_wdata[7:0],io_in_bits_wdata[7:0],io_in_bits_wdata[7:0],
    io_in_bits_wdata[7:0],io_in_bits_wdata[7:0],io_in_bits_wdata[7:0],io_in_bits_wdata[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_92 = {io_in_bits_wdata[15:0],io_in_bits_wdata[15:0],io_in_bits_wdata[15:0],io_in_bits_wdata[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_94 = {io_in_bits_wdata[31:0],io_in_bits_wdata[31:0]}; // @[Cat.scala 30:58]
  wire  _T_95 = 2'h0 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_96 = 2'h1 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_97 = 2'h2 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_98 = 2'h3 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_99 = _T_95 ? _T_89 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_100 = _T_96 ? _T_92 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_101 = _T_97 ? _T_94 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_102 = _T_98 ? io_in_bits_wdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_103 = _T_99 | _T_100; // @[Mux.scala 27:72]
  wire [63:0] _T_104 = _T_103 | _T_101; // @[Mux.scala 27:72]
  wire [1:0] _T_111 = _T_96 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_112 = _T_97 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_113 = _T_98 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_29 = {{1'd0}, _T_95}; // @[Mux.scala 27:72]
  wire [1:0] _T_114 = _GEN_29 | _T_111; // @[Mux.scala 27:72]
  wire [3:0] _GEN_30 = {{2'd0}, _T_114}; // @[Mux.scala 27:72]
  wire [3:0] _T_115 = _GEN_30 | _T_112; // @[Mux.scala 27:72]
  wire [7:0] _GEN_31 = {{4'd0}, _T_115}; // @[Mux.scala 27:72]
  wire [7:0] _T_116 = _GEN_31 | _T_113; // @[Mux.scala 27:72]
  wire [14:0] _GEN_0 = {{7'd0}, _T_116}; // @[SIMD_PipeLSU.scala 92:6]
  wire [14:0] reqWmask = _GEN_0 << exec_addr[2:0]; // @[SIMD_PipeLSU.scala 92:6]
  wire  _T_120 = ~exec_addr[0]; // @[SIMD_PipeLSU.scala 149:32]
  wire  _T_122 = exec_addr[1:0] == 2'h0; // @[SIMD_PipeLSU.scala 150:34]
  wire  _T_124 = exec_addr[2:0] == 3'h0; // @[SIMD_PipeLSU.scala 151:34]
  wire  addrAligned = _T_95 | _T_96 & _T_120 | _T_97 & _T_122 | _T_98 & _T_124; // @[Mux.scala 27:72]
  wire  _T_138 = ~addrAligned; // @[SIMD_PipeLSU.scala 153:57]
  wire  hasloadAddrMisaligned = io_in_valid & _T_28 & ~addrAligned; // @[SIMD_PipeLSU.scala 153:54]
  wire  hasstoreAddrMisaligned = io_in_valid & isStore & _T_138; // @[SIMD_PipeLSU.scala 154:54]
  wire  _T_172 = ~io_dmem_req_bits_cmd[0] & ~io_dmem_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_173 = io_dmem_req_valid & _T_172; // @[SimpleBus.scala 104:29]
  wire  _T_175 = _T_173 & _T_151; // @[SIMD_PipeLSU.scala 175:39]
  reg  hasLoadPF; // @[SIMD_PipeLSU.scala 181:26]
  reg  hasStorePF; // @[SIMD_PipeLSU.scala 182:26]
  wire  _GEN_22 = loadPF_0 & io_in_valid | hasLoadPF; // @[SIMD_PipeLSU.scala 183:30 184:15 181:26]
  wire  _GEN_23 = storePF_0 & io_in_valid | hasStorePF; // @[SIMD_PipeLSU.scala 186:31 187:16 182:26]
  assign io_out_valid = hasLoadPF | hasStorePF | hasloadAddrMisaligned | hasstoreAddrMisaligned | exec_finish; // @[SIMD_PipeLSU.scala 195:83 197:18]
  assign io_out_bits_isMMIO = mmioReg | lsuMMIO_0; // @[SIMD_PipeLSU.scala 79:34]
  assign io_out_bits_loadAddrMisaligned = io_in_valid & _T_28 & ~addrAligned; // @[SIMD_PipeLSU.scala 153:54]
  assign io_out_bits_storeAddrMisaligned = io_in_valid & isStore & _T_138; // @[SIMD_PipeLSU.scala 154:54]
  assign io_out_bits_Decode_cf_pc = io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_exceptionVec_1 = io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_exceptionVec_2 = io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_exceptionVec_12 = io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_0 = io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_1 = io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_2 = io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_3 = io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_4 = io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_5 = io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_6 = io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_7 = io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_8 = io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_9 = io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_10 = io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_intrVec_11 = io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_crossPageIPFFix = io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_cf_runahead_checkpoint_id = io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_ctrl_rfWen = io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_ctrl_rfDest = io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_ctrl_isMou = io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_InstNo = io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_Decode_InstFlag = io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_loadPF = hasLoadPF; // @[SIMD_PipeLSU.scala 193:22]
  assign io_out_bits_storePF = hasStorePF; // @[SIMD_PipeLSU.scala 194:23]
  assign io_out_bits_func = io_in_bits_func; // @[SIMD_PipeLSU.scala 40:15]
  assign io_out_bits_addr = io_in_bits_src1 + io_in_bits_src2; // @[SIMD_PipeLSU.scala 62:26]
  assign io_dmem_req_valid = io_in_valid & req_state == 2'h0 & ~hasloadAddrMisaligned & ~hasstoreAddrMisaligned & ~
    io_flush; // @[SIMD_PipeLSU.scala 161:111]
  assign io_dmem_req_bits_addr = exec_addr[38:0]; // @[SIMD_PipeLSU.scala 144:78]
  assign io_dmem_req_bits_size = {{1'd0}, io_in_bits_func[1:0]}; // @[SimpleBus.scala 66:15]
  assign io_dmem_req_bits_cmd = {{3'd0}, isStore}; // @[SimpleBus.scala 65:14]
  assign io_dmem_req_bits_wmask = reqWmask[7:0]; // @[SimpleBus.scala 68:16]
  assign io_dmem_req_bits_wdata = _T_104 | _T_102; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[SIMD_PipeLSU.scala 124:26]
      req_state <= 2'h0; // @[SIMD_PipeLSU.scala 124:26]
    end else if (io_flush) begin // @[SIMD_PipeLSU.scala 170:17]
      req_state <= 2'h0; // @[SIMD_PipeLSU.scala 170:28]
    end else if (2'h0 == req_state) begin // @[SIMD_PipeLSU.scala 126:22]
      if (_T_40 & ~DTLBPF) begin // @[SIMD_PipeLSU.scala 131:69]
        req_state <= _T_37; // @[SIMD_PipeLSU.scala 131:80]
      end else begin
        req_state <= _GEN_13;
      end
    end else if (2'h1 == req_state) begin // @[SIMD_PipeLSU.scala 126:22]
      req_state <= _GEN_16;
    end else begin
      req_state <= _GEN_18;
    end
    if (reset) begin // @[SIMD_PipeLSU.scala 76:24]
      mmioReg <= 1'h0; // @[SIMD_PipeLSU.scala 76:24]
    end else if (_T) begin // @[SIMD_PipeLSU.scala 78:24]
      mmioReg <= 1'h0; // @[SIMD_PipeLSU.scala 78:34]
    end else if (~mmioReg & io_in_valid) begin // @[SIMD_PipeLSU.scala 77:34]
      mmioReg <= lsuMMIO_0; // @[SIMD_PipeLSU.scala 77:44]
    end
    if (reset) begin // @[SIMD_PipeLSU.scala 181:26]
      hasLoadPF <= 1'h0; // @[SIMD_PipeLSU.scala 181:26]
    end else if (io_flush | _T) begin // @[SIMD_PipeLSU.scala 189:34]
      hasLoadPF <= 1'h0; // @[SIMD_PipeLSU.scala 190:15]
    end else begin
      hasLoadPF <= _GEN_22;
    end
    if (reset) begin // @[SIMD_PipeLSU.scala 182:26]
      hasStorePF <= 1'h0; // @[SIMD_PipeLSU.scala 182:26]
    end else if (io_flush | _T) begin // @[SIMD_PipeLSU.scala 189:34]
      hasStorePF <= 1'h0; // @[SIMD_PipeLSU.scala 191:16]
    end else begin
      hasStorePF <= _GEN_23;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  req_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  mmioReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  hasLoadPF = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  hasStorePF = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_lsu_stage2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_isMMIO,
  input         io_in_bits_loadAddrMisaligned,
  input         io_in_bits_storeAddrMisaligned,
  input  [38:0] io_in_bits_Decode_cf_pc,
  input         io_in_bits_Decode_cf_exceptionVec_1,
  input         io_in_bits_Decode_cf_exceptionVec_2,
  input         io_in_bits_Decode_cf_exceptionVec_12,
  input         io_in_bits_Decode_cf_intrVec_0,
  input         io_in_bits_Decode_cf_intrVec_1,
  input         io_in_bits_Decode_cf_intrVec_2,
  input         io_in_bits_Decode_cf_intrVec_3,
  input         io_in_bits_Decode_cf_intrVec_4,
  input         io_in_bits_Decode_cf_intrVec_5,
  input         io_in_bits_Decode_cf_intrVec_6,
  input         io_in_bits_Decode_cf_intrVec_7,
  input         io_in_bits_Decode_cf_intrVec_8,
  input         io_in_bits_Decode_cf_intrVec_9,
  input         io_in_bits_Decode_cf_intrVec_10,
  input         io_in_bits_Decode_cf_intrVec_11,
  input         io_in_bits_Decode_cf_crossPageIPFFix,
  input  [63:0] io_in_bits_Decode_cf_runahead_checkpoint_id,
  input         io_in_bits_Decode_ctrl_rfWen,
  input  [4:0]  io_in_bits_Decode_ctrl_rfDest,
  input         io_in_bits_Decode_ctrl_isMou,
  input  [4:0]  io_in_bits_Decode_InstNo,
  input         io_in_bits_Decode_InstFlag,
  input         io_in_bits_loadPF,
  input         io_in_bits_storePF,
  input  [6:0]  io_in_bits_func,
  input  [63:0] io_in_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_isMMIO,
  output        io_out_bits_loadAddrMisaligned,
  output        io_out_bits_storeAddrMisaligned,
  output [38:0] io_out_bits_Decode_cf_pc,
  output        io_out_bits_Decode_cf_exceptionVec_1,
  output        io_out_bits_Decode_cf_exceptionVec_2,
  output        io_out_bits_Decode_cf_exceptionVec_12,
  output        io_out_bits_Decode_cf_intrVec_0,
  output        io_out_bits_Decode_cf_intrVec_1,
  output        io_out_bits_Decode_cf_intrVec_2,
  output        io_out_bits_Decode_cf_intrVec_3,
  output        io_out_bits_Decode_cf_intrVec_4,
  output        io_out_bits_Decode_cf_intrVec_5,
  output        io_out_bits_Decode_cf_intrVec_6,
  output        io_out_bits_Decode_cf_intrVec_7,
  output        io_out_bits_Decode_cf_intrVec_8,
  output        io_out_bits_Decode_cf_intrVec_9,
  output        io_out_bits_Decode_cf_intrVec_10,
  output        io_out_bits_Decode_cf_intrVec_11,
  output        io_out_bits_Decode_cf_crossPageIPFFix,
  output [63:0] io_out_bits_Decode_cf_runahead_checkpoint_id,
  output        io_out_bits_Decode_ctrl_rfWen,
  output [4:0]  io_out_bits_Decode_ctrl_rfDest,
  output        io_out_bits_Decode_ctrl_isMou,
  output [4:0]  io_out_bits_Decode_InstNo,
  output        io_out_bits_Decode_InstFlag,
  output        io_out_bits_loadPF,
  output        io_out_bits_storePF,
  output [63:0] io_out_bits_result,
  output [63:0] io_out_bits_addr,
  output        io_dmem_req_valid,
  output [3:0]  io_dmem_req_bits_cmd,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = ~io_in_valid; // @[SIMD_PipeLSU.scala 222:50]
  reg  req_state; // @[SIMD_PipeLSU.scala 245:26]
  wire  _T_146 = io_dmem_resp_ready & io_dmem_resp_valid; // @[Decoupled.scala 40:37]
  wire  exec_finish = req_state | _T_146; // @[SIMD_PipeLSU.scala 295:21]
  wire  _GEN_8 = _T_1 | _T | (_T | ~io_in_valid); // @[SIMD_PipeLSU.scala 222:30 241:{38,51}]
  wire  isStore = io_in_valid & io_in_bits_func[3]; // @[SIMD_PipeLSU.scala 248:28]
  wire  partialLoad = ~isStore & io_in_bits_func != 7'h3; // @[SIMD_PipeLSU.scala 249:30]
  reg [63:0] rdatacache; // @[Reg.scala 15:16]
  wire [63:0] rdataLatch = req_state ? rdatacache : io_dmem_resp_bits_rdata; // @[SIMD_PipeLSU.scala 252:23]
  wire  _T_42 = 3'h0 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_43 = 3'h1 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_44 = 3'h2 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_45 = 3'h3 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_46 = 3'h4 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_47 = 3'h5 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_48 = 3'h6 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_49 = 3'h7 == io_in_bits_addr[2:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_50 = _T_42 ? rdataLatch : 64'h0; // @[Mux.scala 27:72]
  wire [55:0] _T_51 = _T_43 ? rdataLatch[63:8] : 56'h0; // @[Mux.scala 27:72]
  wire [47:0] _T_52 = _T_44 ? rdataLatch[63:16] : 48'h0; // @[Mux.scala 27:72]
  wire [39:0] _T_53 = _T_45 ? rdataLatch[63:24] : 40'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_54 = _T_46 ? rdataLatch[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_55 = _T_47 ? rdataLatch[63:40] : 24'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_56 = _T_48 ? rdataLatch[63:48] : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_57 = _T_49 ? rdataLatch[63:56] : 8'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_21 = {{8'd0}, _T_51}; // @[Mux.scala 27:72]
  wire [63:0] _T_58 = _T_50 | _GEN_21; // @[Mux.scala 27:72]
  wire [63:0] _GEN_22 = {{16'd0}, _T_52}; // @[Mux.scala 27:72]
  wire [63:0] _T_59 = _T_58 | _GEN_22; // @[Mux.scala 27:72]
  wire [63:0] _GEN_23 = {{24'd0}, _T_53}; // @[Mux.scala 27:72]
  wire [63:0] _T_60 = _T_59 | _GEN_23; // @[Mux.scala 27:72]
  wire [63:0] _GEN_24 = {{32'd0}, _T_54}; // @[Mux.scala 27:72]
  wire [63:0] _T_61 = _T_60 | _GEN_24; // @[Mux.scala 27:72]
  wire [63:0] _GEN_25 = {{40'd0}, _T_55}; // @[Mux.scala 27:72]
  wire [63:0] _T_62 = _T_61 | _GEN_25; // @[Mux.scala 27:72]
  wire [63:0] _GEN_26 = {{48'd0}, _T_56}; // @[Mux.scala 27:72]
  wire [63:0] _T_63 = _T_62 | _GEN_26; // @[Mux.scala 27:72]
  wire [63:0] _GEN_27 = {{56'd0}, _T_57}; // @[Mux.scala 27:72]
  wire [63:0] rdataSel = _T_63 | _GEN_27; // @[Mux.scala 27:72]
  wire [55:0] _T_84 = rdataSel[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_85 = {_T_84,rdataSel[7:0]}; // @[Cat.scala 30:58]
  wire [47:0] _T_89 = rdataSel[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_90 = {_T_89,rdataSel[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_94 = rdataSel[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_95 = {_T_94,rdataSel[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_97 = {56'h0,rdataSel[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_99 = {48'h0,rdataSel[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_101 = {32'h0,rdataSel[31:0]}; // @[Cat.scala 30:58]
  wire  _T_102 = 7'h0 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_103 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_104 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_105 = 7'h4 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_106 = 7'h5 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_107 = 7'h6 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_108 = _T_102 ? _T_85 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_109 = _T_103 ? _T_90 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_110 = _T_104 ? _T_95 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_111 = _T_105 ? _T_97 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_112 = _T_106 ? _T_99 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_113 = _T_107 ? _T_101 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_114 = _T_108 | _T_109; // @[Mux.scala 27:72]
  wire [63:0] _T_115 = _T_114 | _T_110; // @[Mux.scala 27:72]
  wire [63:0] _T_116 = _T_115 | _T_111; // @[Mux.scala 27:72]
  wire [63:0] _T_117 = _T_116 | _T_112; // @[Mux.scala 27:72]
  wire [63:0] rdataPartialLoad = _T_117 | _T_113; // @[Mux.scala 27:72]
  wire  _T_139 = exec_finish & io_out_ready; // @[SIMD_PipeLSU.scala 290:79]
  wire  _T_140 = exec_finish & io_out_ready ? 1'h0 : 1'h1; // @[SIMD_PipeLSU.scala 290:66]
  wire  _GEN_11 = _T_139 ? 1'h0 : req_state; // @[SIMD_PipeLSU.scala 245:26 291:{55,66}]
  wire  _T_156 = ~io_dmem_req_bits_cmd[0] & ~io_dmem_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_157 = io_dmem_req_valid & _T_156; // @[SimpleBus.scala 104:29]
  reg  REG_3; // @[StopWatch.scala 24:20]
  wire  _GEN_17 = _T_157 | REG_3; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_160 = io_dmem_req_valid & io_dmem_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  reg  REG_4; // @[StopWatch.scala 24:20]
  wire  _GEN_19 = _T_160 | REG_4; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_163 = io_out_bits_isMMIO & _T; // @[SIMD_PipeLSU.scala 308:44]
  assign io_in_ready = io_in_valid & (io_in_bits_loadPF | io_in_bits_storePF | io_in_bits_loadAddrMisaligned |
    io_in_bits_storeAddrMisaligned) ? 1'h0 : _GEN_8; // @[SIMD_PipeLSU.scala 299:132 301:17]
  assign io_out_valid = io_in_valid & (io_in_bits_loadPF | io_in_bits_storePF | io_in_bits_loadAddrMisaligned |
    io_in_bits_storeAddrMisaligned) | exec_finish; // @[SIMD_PipeLSU.scala 299:132 300:18]
  assign io_out_bits_isMMIO = io_in_bits_isMMIO; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_loadAddrMisaligned = io_in_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_storeAddrMisaligned = io_in_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_pc = io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_exceptionVec_1 = io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_exceptionVec_2 = io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_exceptionVec_12 = io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_0 = io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_1 = io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_2 = io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_3 = io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_4 = io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_5 = io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_6 = io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_7 = io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_8 = io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_9 = io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_10 = io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_intrVec_11 = io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_crossPageIPFFix = io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_cf_runahead_checkpoint_id = io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_ctrl_rfWen = io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_ctrl_rfDest = io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_ctrl_isMou = io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_InstNo = io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_Decode_InstFlag = io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_loadPF = io_in_bits_loadPF; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_storePF = io_in_bits_storePF; // @[SIMD_PipeLSU.scala 214:15]
  assign io_out_bits_result = partialLoad ? rdataPartialLoad : rdataLatch; // @[SIMD_PipeLSU.scala 294:21]
  assign io_out_bits_addr = io_in_bits_addr; // @[SIMD_PipeLSU.scala 214:15]
  assign io_dmem_req_valid = 1'h0;
  assign io_dmem_req_bits_cmd = 4'h0;
  assign io_dmem_resp_ready = 1'h1; // @[SIMD_PipeLSU.scala 297:19]
  always @(posedge clock) begin
    if (reset) begin // @[SIMD_PipeLSU.scala 245:26]
      req_state <= 1'h0; // @[SIMD_PipeLSU.scala 245:26]
    end else if (io_flush) begin // @[SIMD_PipeLSU.scala 304:17]
      req_state <= 1'h0; // @[SIMD_PipeLSU.scala 304:28]
    end else if (~req_state) begin // @[SIMD_PipeLSU.scala 289:22]
      if (_T_146) begin // @[SIMD_PipeLSU.scala 290:48]
        req_state <= _T_140; // @[SIMD_PipeLSU.scala 290:60]
      end
    end else if (req_state) begin // @[SIMD_PipeLSU.scala 289:22]
      req_state <= _GEN_11;
    end
    if (_T_146) begin // @[Reg.scala 16:19]
      rdatacache <= io_dmem_resp_bits_rdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_3 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_146) begin // @[StopWatch.scala 31:19]
      REG_3 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_3 <= _GEN_17;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_4 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_146) begin // @[StopWatch.scala 31:19]
      REG_4 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_4 <= _GEN_19;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  req_state = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  rdatacache = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  REG_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_4 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_lsu_empty_stage(
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_loadAddrMisaligned,
  input         io_in_bits_storeAddrMisaligned,
  input  [38:0] io_in_bits_Decode_cf_pc,
  input         io_in_bits_Decode_cf_exceptionVec_1,
  input         io_in_bits_Decode_cf_exceptionVec_2,
  input         io_in_bits_Decode_cf_exceptionVec_12,
  input         io_in_bits_Decode_cf_intrVec_0,
  input         io_in_bits_Decode_cf_intrVec_1,
  input         io_in_bits_Decode_cf_intrVec_2,
  input         io_in_bits_Decode_cf_intrVec_3,
  input         io_in_bits_Decode_cf_intrVec_4,
  input         io_in_bits_Decode_cf_intrVec_5,
  input         io_in_bits_Decode_cf_intrVec_6,
  input         io_in_bits_Decode_cf_intrVec_7,
  input         io_in_bits_Decode_cf_intrVec_8,
  input         io_in_bits_Decode_cf_intrVec_9,
  input         io_in_bits_Decode_cf_intrVec_10,
  input         io_in_bits_Decode_cf_intrVec_11,
  input         io_in_bits_Decode_cf_crossPageIPFFix,
  input  [63:0] io_in_bits_Decode_cf_runahead_checkpoint_id,
  input         io_in_bits_Decode_ctrl_rfWen,
  input  [4:0]  io_in_bits_Decode_ctrl_rfDest,
  input         io_in_bits_Decode_ctrl_isMou,
  input  [4:0]  io_in_bits_Decode_InstNo,
  input         io_in_bits_Decode_InstFlag,
  input         io_in_bits_loadPF,
  input         io_in_bits_storePF,
  input  [63:0] io_in_bits_result,
  input  [63:0] io_in_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_loadAddrMisaligned,
  output        io_out_bits_storeAddrMisaligned,
  output [38:0] io_out_bits_Decode_cf_pc,
  output        io_out_bits_Decode_cf_exceptionVec_1,
  output        io_out_bits_Decode_cf_exceptionVec_2,
  output        io_out_bits_Decode_cf_exceptionVec_12,
  output        io_out_bits_Decode_cf_intrVec_0,
  output        io_out_bits_Decode_cf_intrVec_1,
  output        io_out_bits_Decode_cf_intrVec_2,
  output        io_out_bits_Decode_cf_intrVec_3,
  output        io_out_bits_Decode_cf_intrVec_4,
  output        io_out_bits_Decode_cf_intrVec_5,
  output        io_out_bits_Decode_cf_intrVec_6,
  output        io_out_bits_Decode_cf_intrVec_7,
  output        io_out_bits_Decode_cf_intrVec_8,
  output        io_out_bits_Decode_cf_intrVec_9,
  output        io_out_bits_Decode_cf_intrVec_10,
  output        io_out_bits_Decode_cf_intrVec_11,
  output        io_out_bits_Decode_cf_crossPageIPFFix,
  output [63:0] io_out_bits_Decode_cf_runahead_checkpoint_id,
  output        io_out_bits_Decode_ctrl_rfWen,
  output [4:0]  io_out_bits_Decode_ctrl_rfDest,
  output        io_out_bits_Decode_ctrl_isMou,
  output [4:0]  io_out_bits_Decode_InstNo,
  output        io_out_bits_Decode_InstFlag,
  output        io_out_bits_loadPF,
  output        io_out_bits_storePF,
  output [63:0] io_out_bits_result,
  output [63:0] io_out_bits_addr
);
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T | ~io_in_valid; // @[SIMD_PipeLSU.scala 313:32]
  assign io_out_valid = io_in_valid; // @[SIMD_PipeLSU.scala 312:16]
  assign io_out_bits_loadAddrMisaligned = io_in_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_storeAddrMisaligned = io_in_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_pc = io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_exceptionVec_1 = io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_exceptionVec_2 = io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_exceptionVec_12 = io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_0 = io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_1 = io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_2 = io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_3 = io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_4 = io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_5 = io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_6 = io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_7 = io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_8 = io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_9 = io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_10 = io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_intrVec_11 = io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_crossPageIPFFix = io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_cf_runahead_checkpoint_id = io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_ctrl_rfWen = io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_ctrl_rfDest = io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_ctrl_isMou = io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_InstNo = io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_Decode_InstFlag = io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_loadPF = io_in_bits_loadPF; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_storePF = io_in_bits_storePF; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_result = io_in_bits_result; // @[SIMD_PipeLSU.scala 314:15]
  assign io_out_bits_addr = io_in_bits_addr; // @[SIMD_PipeLSU.scala 314:15]
endmodule
module AtomALU(
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [6:0]  io_func,
  input         io_isWordOp,
  output [63:0] io_result
);
  wire  isAdderSub = ~io_func[6]; // @[LSU.scala 184:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_src2 ^ _T_2; // @[LSU.scala 185:33]
  wire [64:0] _T_4 = io_src1 + _T_3; // @[LSU.scala 185:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[LSU.scala 185:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[LSU.scala 185:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[LSU.scala 186:21]
  wire  sltu = ~adderRes[64]; // @[LSU.scala 187:14]
  wire  slt = xorRes[63] ^ sltu; // @[LSU.scala 188:28]
  wire [63:0] _T_9 = io_src1 & io_src2; // @[LSU.scala 194:32]
  wire [63:0] _T_10 = io_src1 | io_src2; // @[LSU.scala 195:32]
  wire [63:0] _T_12 = slt ? io_src1 : io_src2; // @[LSU.scala 196:29]
  wire [63:0] _T_14 = slt ? io_src2 : io_src1; // @[LSU.scala 197:29]
  wire [63:0] _T_16 = sltu ? io_src1 : io_src2; // @[LSU.scala 198:29]
  wire [63:0] _T_18 = sltu ? io_src2 : io_src1; // @[LSU.scala 199:29]
  wire [64:0] _T_20 = 6'h22 == io_func[5:0] ? {{1'd0}, io_src2} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_22 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _T_20; // @[Mux.scala 80:57]
  wire [64:0] _T_24 = 6'h25 == io_func[5:0] ? {{1'd0}, _T_9} : _T_22; // @[Mux.scala 80:57]
  wire [64:0] _T_26 = 6'h26 == io_func[5:0] ? {{1'd0}, _T_10} : _T_24; // @[Mux.scala 80:57]
  wire [64:0] _T_28 = 6'h37 == io_func[5:0] ? {{1'd0}, _T_12} : _T_26; // @[Mux.scala 80:57]
  wire [64:0] _T_30 = 6'h30 == io_func[5:0] ? {{1'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire [64:0] _T_32 = 6'h31 == io_func[5:0] ? {{1'd0}, _T_16} : _T_30; // @[Mux.scala 80:57]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _T_18} : _T_32; // @[Mux.scala 80:57]
  wire [31:0] _T_37 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_38 = {_T_37,res[31:0]}; // @[Cat.scala 30:58]
  assign io_result = io_isWordOp ? _T_38 : res[63:0]; // @[LSU.scala 202:20]
endmodule
module lsu_for_atom(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_Decode_cf_instr,
  input  [38:0] io_in_bits_Decode_cf_pc,
  input         io_in_bits_Decode_cf_exceptionVec_1,
  input         io_in_bits_Decode_cf_exceptionVec_2,
  input         io_in_bits_Decode_cf_exceptionVec_12,
  input         io_in_bits_Decode_cf_intrVec_0,
  input         io_in_bits_Decode_cf_intrVec_1,
  input         io_in_bits_Decode_cf_intrVec_2,
  input         io_in_bits_Decode_cf_intrVec_3,
  input         io_in_bits_Decode_cf_intrVec_4,
  input         io_in_bits_Decode_cf_intrVec_5,
  input         io_in_bits_Decode_cf_intrVec_6,
  input         io_in_bits_Decode_cf_intrVec_7,
  input         io_in_bits_Decode_cf_intrVec_8,
  input         io_in_bits_Decode_cf_intrVec_9,
  input         io_in_bits_Decode_cf_intrVec_10,
  input         io_in_bits_Decode_cf_intrVec_11,
  input         io_in_bits_Decode_cf_crossPageIPFFix,
  input  [63:0] io_in_bits_Decode_cf_runahead_checkpoint_id,
  input         io_in_bits_Decode_ctrl_rfWen,
  input  [4:0]  io_in_bits_Decode_ctrl_rfDest,
  input         io_in_bits_Decode_ctrl_isMou,
  input  [4:0]  io_in_bits_Decode_InstNo,
  input         io_in_bits_Decode_InstFlag,
  input  [63:0] io_in_bits_wdata,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_loadAddrMisaligned,
  output        io_out_bits_storeAddrMisaligned,
  output [38:0] io_out_bits_Decode_cf_pc,
  output        io_out_bits_Decode_cf_exceptionVec_1,
  output        io_out_bits_Decode_cf_exceptionVec_2,
  output        io_out_bits_Decode_cf_exceptionVec_12,
  output        io_out_bits_Decode_cf_intrVec_0,
  output        io_out_bits_Decode_cf_intrVec_1,
  output        io_out_bits_Decode_cf_intrVec_2,
  output        io_out_bits_Decode_cf_intrVec_3,
  output        io_out_bits_Decode_cf_intrVec_4,
  output        io_out_bits_Decode_cf_intrVec_5,
  output        io_out_bits_Decode_cf_intrVec_6,
  output        io_out_bits_Decode_cf_intrVec_7,
  output        io_out_bits_Decode_cf_intrVec_8,
  output        io_out_bits_Decode_cf_intrVec_9,
  output        io_out_bits_Decode_cf_intrVec_10,
  output        io_out_bits_Decode_cf_intrVec_11,
  output        io_out_bits_Decode_cf_crossPageIPFFix,
  output [63:0] io_out_bits_Decode_cf_runahead_checkpoint_id,
  output        io_out_bits_Decode_ctrl_rfWen,
  output [4:0]  io_out_bits_Decode_ctrl_rfDest,
  output        io_out_bits_Decode_ctrl_isMou,
  output [4:0]  io_out_bits_Decode_InstNo,
  output        io_out_bits_Decode_InstFlag,
  output        io_out_bits_loadPF,
  output        io_out_bits_storePF,
  output [63:0] io_out_bits_result,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_flush,
  output        setLr_0,
  input         DTLBPF,
  input         loadPF_0,
  input         lr_0,
  output        amoReq_0,
  input         storePF_0,
  input         DTLBENABLE,
  input         DTLBFINISH,
  output [63:0] setLrAddr_0,
  output        setLrVal_0,
  input  [63:0] lr_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] atomALU_io_src1; // @[SIMD_PipeLSU.scala 411:25]
  wire [63:0] atomALU_io_src2; // @[SIMD_PipeLSU.scala 411:25]
  wire [6:0] atomALU_io_func; // @[SIMD_PipeLSU.scala 411:25]
  wire  atomALU_io_isWordOp; // @[SIMD_PipeLSU.scala 411:25]
  wire [63:0] atomALU_io_result; // @[SIMD_PipeLSU.scala 411:25]
  wire  atomReq = io_in_valid & io_in_bits_func[5]; // @[SIMD_PipeLSU.scala 344:26]
  wire  _T_8 = io_in_bits_func == 7'h20; // @[LSU.scala 57:37]
  wire  _T_11 = io_in_bits_func == 7'h21; // @[LSU.scala 58:37]
  wire  _T_13 = io_in_bits_func[5] & ~_T_8 & ~_T_11; // @[LSU.scala 59:61]
  wire  amoReq = io_in_valid & _T_13; // @[SIMD_PipeLSU.scala 345:26]
  wire  lrReq = io_in_valid & _T_8; // @[SIMD_PipeLSU.scala 346:25]
  wire  scReq = io_in_valid & _T_11; // @[SIMD_PipeLSU.scala 347:25]
  wire [2:0] funct3 = io_in_bits_Decode_cf_instr[14:12]; // @[SIMD_PipeLSU.scala 355:44]
  wire  scInvalid = ~(io_in_bits_src1 == lr_addr & lr_0) & scReq; // @[SIMD_PipeLSU.scala 372:46]
  reg  hasLoadPF; // @[SIMD_PipeLSU.scala 388:28]
  reg  hasStorePF; // @[SIMD_PipeLSU.scala 389:28]
  wire  _GEN_0 = loadPF_0 | hasLoadPF; // @[SIMD_PipeLSU.scala 390:17 391:17 388:28]
  wire  _GEN_1 = storePF_0 | hasStorePF; // @[SIMD_PipeLSU.scala 393:18 394:18 389:28]
  wire  _T_27 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [2:0] state; // @[SIMD_PipeLSU.scala 408:24]
  reg [63:0] atomMemReg; // @[SIMD_PipeLSU.scala 409:25]
  reg [63:0] atomRegReg; // @[SIMD_PipeLSU.scala 410:25]
  wire [63:0] _T_36 = io_in_bits_src1 + io_in_bits_src2; // @[SIMD_PipeLSU.scala 423:28]
  reg [1:0] req_state; // @[SIMD_PipeLSU.scala 555:26]
  wire  _T_321 = req_state == 2'h3; // @[SIMD_PipeLSU.scala 623:32]
  wire  _T_322 = io_dmem_resp_ready & io_dmem_resp_valid; // @[Decoupled.scala 40:37]
  wire  exec_finish = req_state == 2'h3 | _T_322 & req_state == 2'h2; // @[SIMD_PipeLSU.scala 623:21]
  wire [2:0] _GEN_4 = amoReq ? 3'h3 : 3'h0; // @[SIMD_PipeLSU.scala 428:15 430:{21,28}]
  wire [2:0] _GEN_5 = lrReq ? 3'h1 : _GEN_4; // @[SIMD_PipeLSU.scala 431:{20,27}]
  wire [2:0] _T_38 = scInvalid ? 3'h0 : 3'h2; // @[SIMD_PipeLSU.scala 432:33]
  wire [1:0] _T_40 = funct3[0] ? 2'h3 : 2'h2; // @[SIMD_PipeLSU.scala 439:26]
  wire [2:0] _GEN_7 = exec_finish ? 3'h4 : state; // @[SIMD_PipeLSU.scala 443:26 444:17 408:24]
  wire [3:0] _T_49 = funct3[0] ? 4'hb : 4'ha; // @[SIMD_PipeLSU.scala 454:26]
  wire [2:0] _GEN_8 = _T_27 ? 3'h0 : state; // @[SIMD_PipeLSU.scala 458:28 459:17 408:24]
  wire [63:0] _GEN_12 = io_in_bits_src1; // @[SIMD_PipeLSU.scala 420:20 477:20]
  wire [6:0] _GEN_13 = 3'h2 == state ? {{3'd0}, _T_49} : io_in_bits_func; // @[SIMD_PipeLSU.scala 420:20 478:20]
  wire  _GEN_15 = 3'h2 == state & io_out_ready; // @[SIMD_PipeLSU.scala 420:20 480:20]
  wire  _GEN_16 = 3'h2 == state & exec_finish; // @[SIMD_PipeLSU.scala 420:20 481:22 417:32]
  wire [2:0] _GEN_17 = 3'h2 == state ? _GEN_8 : state; // @[SIMD_PipeLSU.scala 420:20 408:24]
  wire  _GEN_18 = 3'h1 == state | 3'h2 == state; // @[SIMD_PipeLSU.scala 420:20 464:20]
  wire [6:0] _GEN_20 = 3'h1 == state ? {{5'd0}, _T_40} : _GEN_13; // @[SIMD_PipeLSU.scala 420:20 466:20]
  wire  _GEN_22 = 3'h1 == state ? io_out_ready : _GEN_15; // @[SIMD_PipeLSU.scala 420:20 468:20]
  wire  _GEN_23 = 3'h1 == state ? exec_finish : _GEN_16; // @[SIMD_PipeLSU.scala 420:20 469:22]
  wire [2:0] _GEN_24 = 3'h1 == state ? _GEN_8 : _GEN_17; // @[SIMD_PipeLSU.scala 420:20]
  wire  _GEN_25 = 3'h4 == state | _GEN_18; // @[SIMD_PipeLSU.scala 420:20 452:20]
  wire [6:0] _GEN_27 = 3'h4 == state ? {{3'd0}, _T_49} : _GEN_20; // @[SIMD_PipeLSU.scala 420:20 454:20]
  wire [63:0] _GEN_28 = 3'h4 == state ? atomMemReg : io_in_bits_wdata; // @[SIMD_PipeLSU.scala 420:20 455:20]
  wire  _GEN_29 = 3'h4 == state ? io_out_ready : _GEN_22; // @[SIMD_PipeLSU.scala 420:20 456:20]
  wire  _GEN_30 = 3'h4 == state ? exec_finish : _GEN_23; // @[SIMD_PipeLSU.scala 420:20 457:22]
  wire [2:0] _GEN_31 = 3'h4 == state ? _GEN_8 : _GEN_24; // @[SIMD_PipeLSU.scala 420:20]
  wire  _GEN_32 = 3'h3 == state | _GEN_25; // @[SIMD_PipeLSU.scala 420:20 437:20]
  wire [6:0] _GEN_34 = 3'h3 == state ? {{5'd0}, _T_40} : _GEN_27; // @[SIMD_PipeLSU.scala 420:20 439:20]
  wire [63:0] _GEN_35 = 3'h3 == state ? io_in_bits_wdata : _GEN_28; // @[SIMD_PipeLSU.scala 420:20 440:20]
  wire  _GEN_36 = 3'h3 == state | _GEN_29; // @[SIMD_PipeLSU.scala 420:20 441:20]
  wire  _GEN_37 = 3'h3 == state ? 1'h0 : _GEN_30; // @[SIMD_PipeLSU.scala 420:20 442:22]
  wire  exec_valid = 3'h0 == state ? io_in_valid & ~atomReq : _GEN_32; // @[SIMD_PipeLSU.scala 420:20 422:20]
  wire [6:0] exec_func = 3'h0 == state ? io_in_bits_func : _GEN_34; // @[SIMD_PipeLSU.scala 420:20 424:20]
  wire  isStore = exec_valid & exec_func[3]; // @[SIMD_PipeLSU.scala 551:28]
  wire  _T_116 = ~isStore; // @[SIMD_PipeLSU.scala 552:21]
  wire  partialLoad = ~isStore & exec_func != 7'h3; // @[SIMD_PipeLSU.scala 552:30]
  wire  _T_284 = 7'h0 == exec_func; // @[LookupTree.scala 24:34]
  reg [63:0] addrLatch; // @[SIMD_PipeLSU.scala 550:26]
  wire  _T_224 = 3'h0 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  reg [63:0] rdatacache; // @[Reg.scala 15:16]
  wire [63:0] rdataLatch = _T_321 ? rdatacache : io_dmem_resp_bits_rdata; // @[SIMD_PipeLSU.scala 590:23]
  wire [63:0] _T_232 = _T_224 ? rdataLatch : 64'h0; // @[Mux.scala 27:72]
  wire  _T_225 = 3'h1 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [55:0] _T_233 = _T_225 ? rdataLatch[63:8] : 56'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_70 = {{8'd0}, _T_233}; // @[Mux.scala 27:72]
  wire [63:0] _T_240 = _T_232 | _GEN_70; // @[Mux.scala 27:72]
  wire  _T_226 = 3'h2 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [47:0] _T_234 = _T_226 ? rdataLatch[63:16] : 48'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_71 = {{16'd0}, _T_234}; // @[Mux.scala 27:72]
  wire [63:0] _T_241 = _T_240 | _GEN_71; // @[Mux.scala 27:72]
  wire  _T_227 = 3'h3 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [39:0] _T_235 = _T_227 ? rdataLatch[63:24] : 40'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_72 = {{24'd0}, _T_235}; // @[Mux.scala 27:72]
  wire [63:0] _T_242 = _T_241 | _GEN_72; // @[Mux.scala 27:72]
  wire  _T_228 = 3'h4 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_236 = _T_228 ? rdataLatch[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_73 = {{32'd0}, _T_236}; // @[Mux.scala 27:72]
  wire [63:0] _T_243 = _T_242 | _GEN_73; // @[Mux.scala 27:72]
  wire  _T_229 = 3'h5 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [23:0] _T_237 = _T_229 ? rdataLatch[63:40] : 24'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_74 = {{40'd0}, _T_237}; // @[Mux.scala 27:72]
  wire [63:0] _T_244 = _T_243 | _GEN_74; // @[Mux.scala 27:72]
  wire  _T_230 = 3'h6 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [15:0] _T_238 = _T_230 ? rdataLatch[63:48] : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_75 = {{48'd0}, _T_238}; // @[Mux.scala 27:72]
  wire [63:0] _T_245 = _T_244 | _GEN_75; // @[Mux.scala 27:72]
  wire  _T_231 = 3'h7 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [7:0] _T_239 = _T_231 ? rdataLatch[63:56] : 8'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_76 = {{56'd0}, _T_239}; // @[Mux.scala 27:72]
  wire [63:0] rdataSel = _T_245 | _GEN_76; // @[Mux.scala 27:72]
  wire [55:0] _T_266 = rdataSel[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_267 = {_T_266,rdataSel[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_290 = _T_284 ? _T_267 : 64'h0; // @[Mux.scala 27:72]
  wire  _T_285 = 7'h1 == exec_func; // @[LookupTree.scala 24:34]
  wire [47:0] _T_271 = rdataSel[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_272 = {_T_271,rdataSel[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_291 = _T_285 ? _T_272 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_296 = _T_290 | _T_291; // @[Mux.scala 27:72]
  wire  _T_286 = 7'h2 == exec_func; // @[LookupTree.scala 24:34]
  wire [31:0] _T_276 = rdataSel[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_277 = {_T_276,rdataSel[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_292 = _T_286 ? _T_277 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_297 = _T_296 | _T_292; // @[Mux.scala 27:72]
  wire  _T_287 = 7'h4 == exec_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_279 = {56'h0,rdataSel[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_293 = _T_287 ? _T_279 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_298 = _T_297 | _T_293; // @[Mux.scala 27:72]
  wire  _T_288 = 7'h5 == exec_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_281 = {48'h0,rdataSel[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_294 = _T_288 ? _T_281 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_299 = _T_298 | _T_294; // @[Mux.scala 27:72]
  wire  _T_289 = 7'h6 == exec_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_283 = {32'h0,rdataSel[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_295 = _T_289 ? _T_283 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] rdataPartialLoad = _T_299 | _T_295; // @[Mux.scala 27:72]
  wire [63:0] exec_result = partialLoad ? rdataPartialLoad : rdataLatch; // @[SIMD_PipeLSU.scala 622:21]
  wire [63:0] exec_addr = 3'h0 == state ? _T_36 : io_in_bits_src1; // @[SIMD_PipeLSU.scala 420:20 423:20]
  wire [63:0] exec_wdata = 3'h0 == state ? io_in_bits_wdata : _GEN_35; // @[SIMD_PipeLSU.scala 420:20 425:20]
  wire  exec_clear = 3'h0 == state ? io_out_ready : _GEN_36; // @[SIMD_PipeLSU.scala 420:20 426:20]
  wire  _GEN_46 = 3'h0 == state ? exec_finish | scInvalid : _GEN_37; // @[SIMD_PipeLSU.scala 420:20 427:23]
  wire [63:0] _T_101 = state == 3'h4 ? atomRegReg : exec_result; // @[SIMD_PipeLSU.scala 502:52]
  wire  _T_119 = io_dmem_req_ready & io_dmem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_120 = _T_119 & DTLBENABLE; // @[SIMD_PipeLSU.scala 559:29]
  wire [1:0] _GEN_56 = _T_119 & DTLBENABLE ? 2'h1 : req_state; // @[SIMD_PipeLSU.scala 555:26 559:{45,57}]
  wire [1:0] _GEN_57 = _T_119 & ~DTLBENABLE ? 2'h2 : _GEN_56; // @[SIMD_PipeLSU.scala 560:{45,57}]
  wire  _T_126 = _T_120 & DTLBFINISH; // @[SIMD_PipeLSU.scala 561:43]
  wire [1:0] _GEN_58 = _T_120 & DTLBFINISH & DTLBPF ? 2'h0 : _GEN_57; // @[SIMD_PipeLSU.scala 561:{68,79}]
  wire  _T_131 = ~DTLBPF; // @[SIMD_PipeLSU.scala 562:60]
  wire [1:0] _GEN_60 = DTLBFINISH & DTLBPF ? 2'h0 : req_state; // @[SIMD_PipeLSU.scala 555:26 565:{36,48}]
  wire [1:0] _GEN_61 = DTLBFINISH & _T_131 ? 2'h2 : _GEN_60; // @[SIMD_PipeLSU.scala 566:{36,48}]
  wire  _T_139 = exec_finish & exec_clear; // @[SIMD_PipeLSU.scala 568:79]
  wire [1:0] _T_140 = exec_finish & exec_clear ? 2'h0 : 2'h3; // @[SIMD_PipeLSU.scala 568:66]
  wire [1:0] _GEN_62 = _T_322 ? _T_140 : req_state; // @[SIMD_PipeLSU.scala 555:26 568:{48,60}]
  wire [1:0] _GEN_63 = _T_139 ? 2'h0 : req_state; // @[SIMD_PipeLSU.scala 555:26 569:{55,66}]
  wire [1:0] _GEN_64 = 2'h3 == req_state ? _GEN_63 : req_state; // @[SIMD_PipeLSU.scala 557:22 555:26]
  wire [1:0] _GEN_65 = 2'h2 == req_state ? _GEN_62 : _GEN_64; // @[SIMD_PipeLSU.scala 557:22]
  wire [63:0] _T_175 = {exec_wdata[7:0],exec_wdata[7:0],exec_wdata[7:0],exec_wdata[7:0],exec_wdata[7:0],exec_wdata[7:0],
    exec_wdata[7:0],exec_wdata[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_178 = {exec_wdata[15:0],exec_wdata[15:0],exec_wdata[15:0],exec_wdata[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_180 = {exec_wdata[31:0],exec_wdata[31:0]}; // @[Cat.scala 30:58]
  wire  _T_181 = 2'h0 == exec_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_182 = 2'h1 == exec_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_183 = 2'h2 == exec_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_184 = 2'h3 == exec_func[1:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_185 = _T_181 ? _T_175 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_186 = _T_182 ? _T_178 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_187 = _T_183 ? _T_180 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_188 = _T_184 ? exec_wdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_189 = _T_185 | _T_186; // @[Mux.scala 27:72]
  wire [63:0] _T_190 = _T_189 | _T_187; // @[Mux.scala 27:72]
  wire [1:0] _T_197 = _T_182 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_198 = _T_183 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_199 = _T_184 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_77 = {{1'd0}, _T_181}; // @[Mux.scala 27:72]
  wire [1:0] _T_200 = _GEN_77 | _T_197; // @[Mux.scala 27:72]
  wire [3:0] _GEN_78 = {{2'd0}, _T_200}; // @[Mux.scala 27:72]
  wire [3:0] _T_201 = _GEN_78 | _T_198; // @[Mux.scala 27:72]
  wire [7:0] _GEN_79 = {{4'd0}, _T_201}; // @[Mux.scala 27:72]
  wire [7:0] _T_202 = _GEN_79 | _T_199; // @[Mux.scala 27:72]
  wire [14:0] _GEN_9 = {{7'd0}, _T_202}; // @[SIMD_PipeLSU.scala 523:8]
  wire [14:0] reqWmask = _GEN_9 << exec_addr[2:0]; // @[SIMD_PipeLSU.scala 523:8]
  wire  _T_303 = ~exec_addr[0]; // @[SIMD_PipeLSU.scala 618:32]
  wire  _T_305 = exec_addr[1:0] == 2'h0; // @[SIMD_PipeLSU.scala 619:34]
  wire  _T_307 = exec_addr[2:0] == 3'h0; // @[SIMD_PipeLSU.scala 620:34]
  wire  addrAligned = _T_181 | _T_182 & _T_303 | _T_183 & _T_305 | _T_184 & _T_307; // @[Mux.scala 27:72]
  wire  _T_337 = ~addrAligned; // @[SIMD_PipeLSU.scala 629:74]
  wire  setLr = _T_27 & (lrReq | scReq); // @[SIMD_PipeLSU.scala 498:28]
  wire  setLrVal = lrReq; // @[SIMD_PipeLSU.scala 346:25]
  wire [63:0] setLrAddr = io_in_bits_src1; // @[SIMD_PipeLSU.scala 363:25 500:15]
  AtomALU atomALU ( // @[SIMD_PipeLSU.scala 411:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io_out_valid = io_in_valid & (io_out_bits_storePF | io_out_bits_loadPF | io_out_bits_loadAddrMisaligned |
    io_out_bits_storeAddrMisaligned) | _GEN_46; // @[SIMD_PipeLSU.scala 488:138 490:20]
  assign io_out_bits_loadAddrMisaligned = exec_valid & _T_116 & ~amoReq & ~addrAligned; // @[SIMD_PipeLSU.scala 629:71]
  assign io_out_bits_storeAddrMisaligned = exec_valid & (isStore | amoReq) & _T_337; // @[SIMD_PipeLSU.scala 630:71]
  assign io_out_bits_Decode_cf_pc = io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_exceptionVec_1 = io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_exceptionVec_2 = io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_exceptionVec_12 = io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_0 = io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_1 = io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_2 = io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_3 = io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_4 = io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_5 = io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_6 = io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_7 = io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_8 = io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_9 = io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_10 = io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_intrVec_11 = io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_crossPageIPFFix = io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_cf_runahead_checkpoint_id = io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_ctrl_rfWen = io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_ctrl_rfDest = io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_ctrl_isMou = io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_InstNo = io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_Decode_InstFlag = io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 340:17]
  assign io_out_bits_loadPF = hasLoadPF; // @[SIMD_PipeLSU.scala 400:24]
  assign io_out_bits_storePF = hasStorePF; // @[SIMD_PipeLSU.scala 401:25]
  assign io_out_bits_result = scReq ? {{63'd0}, scInvalid} : _T_101; // @[SIMD_PipeLSU.scala 502:30]
  assign io_dmem_req_valid = exec_valid & req_state == 2'h0 & ~io_out_bits_loadAddrMisaligned & ~
    io_out_bits_storeAddrMisaligned & ~io_flush; // @[SIMD_PipeLSU.scala 585:129]
  assign io_dmem_req_bits_addr = exec_addr[38:0]; // @[SIMD_PipeLSU.scala 576:78]
  assign io_dmem_req_bits_size = {{1'd0}, exec_func[1:0]}; // @[SimpleBus.scala 66:15]
  assign io_dmem_req_bits_cmd = {{3'd0}, isStore}; // @[SimpleBus.scala 65:14]
  assign io_dmem_req_bits_wmask = reqWmask[7:0]; // @[SimpleBus.scala 68:16]
  assign io_dmem_req_bits_wdata = _T_190 | _T_188; // @[Mux.scala 27:72]
  assign io_dmem_resp_ready = 1'h1; // @[SIMD_PipeLSU.scala 586:19]
  assign setLr_0 = setLr;
  assign amoReq_0 = amoReq;
  assign setLrAddr_0 = _GEN_12;
  assign setLrVal_0 = setLrVal;
  assign atomALU_io_src1 = partialLoad ? rdataPartialLoad : rdataLatch; // @[SIMD_PipeLSU.scala 622:21]
  assign atomALU_io_src2 = io_in_bits_wdata; // @[SIMD_PipeLSU.scala 413:21]
  assign atomALU_io_func = io_in_bits_func; // @[SIMD_PipeLSU.scala 414:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[SIMD_PipeLSU.scala 357:22]
  always @(posedge clock) begin
    if (reset) begin // @[SIMD_PipeLSU.scala 388:28]
      hasLoadPF <= 1'h0; // @[SIMD_PipeLSU.scala 388:28]
    end else if (io_flush | _T_27) begin // @[SIMD_PipeLSU.scala 396:36]
      hasLoadPF <= 1'h0; // @[SIMD_PipeLSU.scala 397:17]
    end else begin
      hasLoadPF <= _GEN_0;
    end
    if (reset) begin // @[SIMD_PipeLSU.scala 389:28]
      hasStorePF <= 1'h0; // @[SIMD_PipeLSU.scala 389:28]
    end else if (io_flush | _T_27) begin // @[SIMD_PipeLSU.scala 396:36]
      hasStorePF <= 1'h0; // @[SIMD_PipeLSU.scala 398:18]
    end else begin
      hasStorePF <= _GEN_1;
    end
    if (reset) begin // @[SIMD_PipeLSU.scala 408:24]
      state <= 3'h0; // @[SIMD_PipeLSU.scala 408:24]
    end else if (io_flush) begin // @[SIMD_PipeLSU.scala 514:19]
      state <= 3'h0; // @[SIMD_PipeLSU.scala 514:26]
    end else if (3'h0 == state) begin // @[SIMD_PipeLSU.scala 420:20]
      if (scReq) begin // @[SIMD_PipeLSU.scala 432:20]
        state <= _T_38; // @[SIMD_PipeLSU.scala 432:27]
      end else begin
        state <= _GEN_5;
      end
    end else if (3'h3 == state) begin // @[SIMD_PipeLSU.scala 420:20]
      state <= _GEN_7;
    end else begin
      state <= _GEN_31;
    end
    if (!(3'h0 == state)) begin // @[SIMD_PipeLSU.scala 420:20]
      if (3'h3 == state) begin // @[SIMD_PipeLSU.scala 420:20]
        atomMemReg <= atomALU_io_result; // @[SIMD_PipeLSU.scala 447:20]
      end
    end
    if (!(3'h0 == state)) begin // @[SIMD_PipeLSU.scala 420:20]
      if (3'h3 == state) begin // @[SIMD_PipeLSU.scala 420:20]
        if (partialLoad) begin // @[SIMD_PipeLSU.scala 622:21]
          atomRegReg <= rdataPartialLoad;
        end else if (_T_321) begin // @[SIMD_PipeLSU.scala 590:23]
          atomRegReg <= rdatacache;
        end else begin
          atomRegReg <= io_dmem_resp_bits_rdata;
        end
      end
    end
    if (reset) begin // @[SIMD_PipeLSU.scala 555:26]
      req_state <= 2'h0; // @[SIMD_PipeLSU.scala 555:26]
    end else if (io_flush) begin // @[SIMD_PipeLSU.scala 632:17]
      req_state <= 2'h0; // @[SIMD_PipeLSU.scala 632:28]
    end else if (2'h0 == req_state) begin // @[SIMD_PipeLSU.scala 557:22]
      if (_T_126 & ~DTLBPF) begin // @[SIMD_PipeLSU.scala 562:69]
        req_state <= 2'h2; // @[SIMD_PipeLSU.scala 562:80]
      end else begin
        req_state <= _GEN_58;
      end
    end else if (2'h1 == req_state) begin // @[SIMD_PipeLSU.scala 557:22]
      req_state <= _GEN_61;
    end else begin
      req_state <= _GEN_65;
    end
    if (3'h0 == state) begin // @[SIMD_PipeLSU.scala 420:20]
      addrLatch <= _T_36; // @[SIMD_PipeLSU.scala 423:20]
    end else begin
      addrLatch <= io_in_bits_src1;
    end
    if (_T_322) begin // @[Reg.scala 16:19]
      rdatacache <= io_dmem_resp_bits_rdata; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasLoadPF = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hasStorePF = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  atomMemReg = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  atomRegReg = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  req_state = _RAND_5[1:0];
  _RAND_6 = {2{`RANDOM}};
  addrLatch = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rdatacache = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_lsu_atom(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_wdata,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  output        io_loadAddrMisaligned,
  output        io_storeAddrMisaligned,
  input         io_flush,
  output [38:0] io_DecodeOut_cf_pc,
  output        io_DecodeOut_cf_exceptionVec_1,
  output        io_DecodeOut_cf_exceptionVec_2,
  output        io_DecodeOut_cf_exceptionVec_12,
  output        io_DecodeOut_cf_intrVec_0,
  output        io_DecodeOut_cf_intrVec_1,
  output        io_DecodeOut_cf_intrVec_2,
  output        io_DecodeOut_cf_intrVec_3,
  output        io_DecodeOut_cf_intrVec_4,
  output        io_DecodeOut_cf_intrVec_5,
  output        io_DecodeOut_cf_intrVec_6,
  output        io_DecodeOut_cf_intrVec_7,
  output        io_DecodeOut_cf_intrVec_8,
  output        io_DecodeOut_cf_intrVec_9,
  output        io_DecodeOut_cf_intrVec_10,
  output        io_DecodeOut_cf_intrVec_11,
  output        io_DecodeOut_cf_crossPageIPFFix,
  output [63:0] io_DecodeOut_cf_runahead_checkpoint_id,
  output        io_DecodeOut_ctrl_rfWen,
  output [4:0]  io_DecodeOut_ctrl_rfDest,
  output        io_DecodeOut_ctrl_isMou,
  output [4:0]  io_DecodeOut_InstNo,
  output        io_DecodeOut_InstFlag,
  input  [63:0] io_DecodeIn_cf_instr,
  input  [38:0] io_DecodeIn_cf_pc,
  input         io_DecodeIn_cf_exceptionVec_1,
  input         io_DecodeIn_cf_exceptionVec_2,
  input         io_DecodeIn_cf_exceptionVec_12,
  input         io_DecodeIn_cf_intrVec_0,
  input         io_DecodeIn_cf_intrVec_1,
  input         io_DecodeIn_cf_intrVec_2,
  input         io_DecodeIn_cf_intrVec_3,
  input         io_DecodeIn_cf_intrVec_4,
  input         io_DecodeIn_cf_intrVec_5,
  input         io_DecodeIn_cf_intrVec_6,
  input         io_DecodeIn_cf_intrVec_7,
  input         io_DecodeIn_cf_intrVec_8,
  input         io_DecodeIn_cf_intrVec_9,
  input         io_DecodeIn_cf_intrVec_10,
  input         io_DecodeIn_cf_intrVec_11,
  input         io_DecodeIn_cf_crossPageIPFFix,
  input  [63:0] io_DecodeIn_cf_runahead_checkpoint_id,
  input         io_DecodeIn_ctrl_rfWen,
  input  [4:0]  io_DecodeIn_ctrl_rfDest,
  input         io_DecodeIn_ctrl_isMou,
  input  [4:0]  io_DecodeIn_InstNo,
  input         io_DecodeIn_InstFlag,
  output        io_loadPF,
  output        io_storePF,
  output        lsu_firststage_fire_0,
  output        setLr,
  input         _T_408,
  input         io_memMMU_dmem_loadPF,
  input         ismmio,
  input         lr,
  output        amoReq,
  input         io_memMMU_dmem_storePF,
  input         vmEnable,
  output [63:0] addr_0,
  input         _T_407,
  output [63:0] setLrAddr,
  output        setLrVal,
  input  [63:0] lrAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
`endif // RANDOMIZE_REG_INIT
  wire  stage1_clock; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_reset; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_valid; // @[SIMD_PipeLSU.scala 652:22]
  wire [38:0] stage1_io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 652:22]
  wire [4:0] stage1_io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 652:22]
  wire [4:0] stage1_io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_in_bits_wdata; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_in_bits_src1; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_in_bits_src2; // @[SIMD_PipeLSU.scala 652:22]
  wire [6:0] stage1_io_in_bits_func; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_ready; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_valid; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_isMMIO; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 652:22]
  wire [38:0] stage1_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 652:22]
  wire [4:0] stage1_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 652:22]
  wire [4:0] stage1_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 652:22]
  wire [6:0] stage1_io_out_bits_func; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_out_bits_addr; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_dmem_req_ready; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_dmem_req_valid; // @[SIMD_PipeLSU.scala 652:22]
  wire [38:0] stage1_io_dmem_req_bits_addr; // @[SIMD_PipeLSU.scala 652:22]
  wire [2:0] stage1_io_dmem_req_bits_size; // @[SIMD_PipeLSU.scala 652:22]
  wire [3:0] stage1_io_dmem_req_bits_cmd; // @[SIMD_PipeLSU.scala 652:22]
  wire [7:0] stage1_io_dmem_req_bits_wmask; // @[SIMD_PipeLSU.scala 652:22]
  wire [63:0] stage1_io_dmem_req_bits_wdata; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_io_flush; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_DTLBPF; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_loadPF_0; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_lsuMMIO_0; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_storePF_0; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_DTLBENABLE; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage1_DTLBFINISH; // @[SIMD_PipeLSU.scala 652:22]
  wire  stage2_clock; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_reset; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_ready; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_valid; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_isMMIO; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 653:22]
  wire [38:0] stage2_io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 653:22]
  wire [63:0] stage2_io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 653:22]
  wire [4:0] stage2_io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 653:22]
  wire [4:0] stage2_io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_loadPF; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_in_bits_storePF; // @[SIMD_PipeLSU.scala 653:22]
  wire [6:0] stage2_io_in_bits_func; // @[SIMD_PipeLSU.scala 653:22]
  wire [63:0] stage2_io_in_bits_addr; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_ready; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_valid; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_isMMIO; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 653:22]
  wire [38:0] stage2_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 653:22]
  wire [63:0] stage2_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 653:22]
  wire [4:0] stage2_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 653:22]
  wire [4:0] stage2_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 653:22]
  wire [63:0] stage2_io_out_bits_result; // @[SIMD_PipeLSU.scala 653:22]
  wire [63:0] stage2_io_out_bits_addr; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_dmem_req_valid; // @[SIMD_PipeLSU.scala 653:22]
  wire [3:0] stage2_io_dmem_req_bits_cmd; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_dmem_resp_ready; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_dmem_resp_valid; // @[SIMD_PipeLSU.scala 653:22]
  wire [63:0] stage2_io_dmem_resp_bits_rdata; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage2_io_flush; // @[SIMD_PipeLSU.scala 653:22]
  wire  stage_empty_io_in_ready; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_valid; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 654:27]
  wire [38:0] stage_empty_io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 654:27]
  wire [63:0] stage_empty_io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 654:27]
  wire [4:0] stage_empty_io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 654:27]
  wire [4:0] stage_empty_io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_loadPF; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_in_bits_storePF; // @[SIMD_PipeLSU.scala 654:27]
  wire [63:0] stage_empty_io_in_bits_result; // @[SIMD_PipeLSU.scala 654:27]
  wire [63:0] stage_empty_io_in_bits_addr; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_ready; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_valid; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 654:27]
  wire [38:0] stage_empty_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 654:27]
  wire [63:0] stage_empty_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 654:27]
  wire [4:0] stage_empty_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 654:27]
  wire [4:0] stage_empty_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 654:27]
  wire  stage_empty_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 654:27]
  wire [63:0] stage_empty_io_out_bits_result; // @[SIMD_PipeLSU.scala 654:27]
  wire [63:0] stage_empty_io_out_bits_addr; // @[SIMD_PipeLSU.scala 654:27]
  wire  atomstage_clock; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_reset; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_valid; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_in_bits_Decode_cf_instr; // @[SIMD_PipeLSU.scala 655:25]
  wire [38:0] atomstage_io_in_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_in_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 655:25]
  wire [4:0] atomstage_io_in_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 655:25]
  wire [4:0] atomstage_io_in_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_in_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_in_bits_wdata; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_in_bits_src1; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_in_bits_src2; // @[SIMD_PipeLSU.scala 655:25]
  wire [6:0] atomstage_io_in_bits_func; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_ready; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_valid; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 655:25]
  wire [38:0] atomstage_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 655:25]
  wire [4:0] atomstage_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 655:25]
  wire [4:0] atomstage_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_out_bits_result; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_dmem_req_ready; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_dmem_req_valid; // @[SIMD_PipeLSU.scala 655:25]
  wire [38:0] atomstage_io_dmem_req_bits_addr; // @[SIMD_PipeLSU.scala 655:25]
  wire [2:0] atomstage_io_dmem_req_bits_size; // @[SIMD_PipeLSU.scala 655:25]
  wire [3:0] atomstage_io_dmem_req_bits_cmd; // @[SIMD_PipeLSU.scala 655:25]
  wire [7:0] atomstage_io_dmem_req_bits_wmask; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_dmem_req_bits_wdata; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_dmem_resp_ready; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_dmem_resp_valid; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_io_dmem_resp_bits_rdata; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_io_flush; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_setLr_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_DTLBPF; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_loadPF_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_lr_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_amoReq_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_storePF_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_DTLBENABLE; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_DTLBFINISH; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_setLrAddr_0; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomstage_setLrVal_0; // @[SIMD_PipeLSU.scala 655:25]
  wire [63:0] atomstage_lr_addr; // @[SIMD_PipeLSU.scala 655:25]
  wire  atomReq = io_in_bits_func[5]; // @[LSU.scala 54:38]
  wire  stage2_exp = stage2_io_in_valid & (stage2_io_out_bits_loadAddrMisaligned |
    stage2_io_out_bits_storeAddrMisaligned | stage2_io_out_bits_storePF | stage2_io_out_bits_loadPF); // @[SIMD_PipeLSU.scala 687:37]
  wire  _T = ~stage2_exp; // @[SIMD_PipeLSU.scala 667:34]
  wire  stage_empty_exp = stage_empty_io_in_valid & (stage_empty_io_out_bits_loadAddrMisaligned |
    stage_empty_io_out_bits_storeAddrMisaligned | stage_empty_io_out_bits_storePF | stage_empty_io_out_bits_loadPF); // @[SIMD_PipeLSU.scala 691:46]
  wire  _T_6 = stage2_io_in_valid ? stage2_io_out_ready : 1'h1; // @[SIMD_PipeLSU.scala 667:84]
  wire  _T_11 = stage2_io_out_ready & stage2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_11 ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_12 = stage1_io_out_valid & stage2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = stage1_io_out_valid & stage2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg  r_isMMIO; // @[Reg.scala 15:16]
  reg  r_loadAddrMisaligned; // @[Reg.scala 15:16]
  reg  r_storeAddrMisaligned; // @[Reg.scala 15:16]
  reg [38:0] r_Decode_cf_pc; // @[Reg.scala 15:16]
  reg  r_Decode_cf_exceptionVec_1; // @[Reg.scala 15:16]
  reg  r_Decode_cf_exceptionVec_2; // @[Reg.scala 15:16]
  reg  r_Decode_cf_exceptionVec_12; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_0; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_1; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_2; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_3; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_4; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_5; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_6; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_7; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_8; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_9; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_10; // @[Reg.scala 15:16]
  reg  r_Decode_cf_intrVec_11; // @[Reg.scala 15:16]
  reg  r_Decode_cf_crossPageIPFFix; // @[Reg.scala 15:16]
  reg [63:0] r_Decode_cf_runahead_checkpoint_id; // @[Reg.scala 15:16]
  reg  r_Decode_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] r_Decode_ctrl_rfDest; // @[Reg.scala 15:16]
  reg  r_Decode_ctrl_isMou; // @[Reg.scala 15:16]
  reg [4:0] r_Decode_InstNo; // @[Reg.scala 15:16]
  reg  r_Decode_InstFlag; // @[Reg.scala 15:16]
  reg  r_loadPF; // @[Reg.scala 15:16]
  reg  r_storePF; // @[Reg.scala 15:16]
  reg [6:0] r_func; // @[Reg.scala 15:16]
  reg [63:0] r_addr; // @[Reg.scala 15:16]
  wire  _GEN_80 = stage2_io_in_valid & stage2_exp & stage2_io_out_valid; // @[SIMD_PipeLSU.scala 707:47 708:21]
  wire  _GEN_87 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_88 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_89 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_96 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_104 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_118 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_121 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_122 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_123 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_124 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_125 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_126 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_127 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_128 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_129 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_130 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_131 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_132 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_134 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_135 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_145 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_155 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  _GEN_156 = stage2_io_in_valid & stage2_exp & stage2_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 707:47 709:21]
  wire  empty_out_ready = stage_empty_io_in_ready;
  wire  _GEN_158 = stage2_io_in_valid & stage2_exp ? empty_out_ready : io_out_ready; // @[SIMD_PipeLSU.scala 689:23 707:47 710:25]
  wire  empty_out_valid = atomstage_io_in_valid ? atomstage_io_out_valid : _GEN_80; // @[SIMD_PipeLSU.scala 703:30 704:21]
  wire  _T_23 = stage_empty_io_out_ready & stage_empty_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_239 = _T_23 ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_24 = empty_out_valid & stage_empty_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_240 = empty_out_valid & stage_empty_io_in_ready | _GEN_239; // @[Pipeline.scala 26:{38,46}]
  reg  r_1_loadAddrMisaligned; // @[Reg.scala 15:16]
  reg  r_1_storeAddrMisaligned; // @[Reg.scala 15:16]
  reg [38:0] r_1_Decode_cf_pc; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_exceptionVec_1; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_exceptionVec_2; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_exceptionVec_12; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_0; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_1; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_2; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_3; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_4; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_5; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_6; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_7; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_8; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_9; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_10; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_intrVec_11; // @[Reg.scala 15:16]
  reg  r_1_Decode_cf_crossPageIPFFix; // @[Reg.scala 15:16]
  reg [63:0] r_1_Decode_cf_runahead_checkpoint_id; // @[Reg.scala 15:16]
  reg  r_1_Decode_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] r_1_Decode_ctrl_rfDest; // @[Reg.scala 15:16]
  reg  r_1_Decode_ctrl_isMou; // @[Reg.scala 15:16]
  reg [4:0] r_1_Decode_InstNo; // @[Reg.scala 15:16]
  reg  r_1_Decode_InstFlag; // @[Reg.scala 15:16]
  reg  r_1_loadPF; // @[Reg.scala 15:16]
  reg  r_1_storePF; // @[Reg.scala 15:16]
  reg [63:0] r_1_result; // @[Reg.scala 15:16]
  reg [63:0] r_1_addr; // @[Reg.scala 15:16]
  wire  _T_32 = atomstage_io_out_ready & atomstage_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = stage1_io_out_ready & stage1_io_out_valid; // @[Decoupled.scala 40:37]
  wire  lsu_firststage_fire = atomstage_io_in_valid ? _T_32 : _T_33; // @[SIMD_PipeLSU.scala 731:30 733:25 739:25]
  wire [63:0] addr = stage_empty_io_out_bits_addr;
  pipeline_lsu_stage1 stage1 ( // @[SIMD_PipeLSU.scala 652:22]
    .clock(stage1_clock),
    .reset(stage1_reset),
    .io_in_valid(stage1_io_in_valid),
    .io_in_bits_Decode_cf_pc(stage1_io_in_bits_Decode_cf_pc),
    .io_in_bits_Decode_cf_exceptionVec_1(stage1_io_in_bits_Decode_cf_exceptionVec_1),
    .io_in_bits_Decode_cf_exceptionVec_2(stage1_io_in_bits_Decode_cf_exceptionVec_2),
    .io_in_bits_Decode_cf_exceptionVec_12(stage1_io_in_bits_Decode_cf_exceptionVec_12),
    .io_in_bits_Decode_cf_intrVec_0(stage1_io_in_bits_Decode_cf_intrVec_0),
    .io_in_bits_Decode_cf_intrVec_1(stage1_io_in_bits_Decode_cf_intrVec_1),
    .io_in_bits_Decode_cf_intrVec_2(stage1_io_in_bits_Decode_cf_intrVec_2),
    .io_in_bits_Decode_cf_intrVec_3(stage1_io_in_bits_Decode_cf_intrVec_3),
    .io_in_bits_Decode_cf_intrVec_4(stage1_io_in_bits_Decode_cf_intrVec_4),
    .io_in_bits_Decode_cf_intrVec_5(stage1_io_in_bits_Decode_cf_intrVec_5),
    .io_in_bits_Decode_cf_intrVec_6(stage1_io_in_bits_Decode_cf_intrVec_6),
    .io_in_bits_Decode_cf_intrVec_7(stage1_io_in_bits_Decode_cf_intrVec_7),
    .io_in_bits_Decode_cf_intrVec_8(stage1_io_in_bits_Decode_cf_intrVec_8),
    .io_in_bits_Decode_cf_intrVec_9(stage1_io_in_bits_Decode_cf_intrVec_9),
    .io_in_bits_Decode_cf_intrVec_10(stage1_io_in_bits_Decode_cf_intrVec_10),
    .io_in_bits_Decode_cf_intrVec_11(stage1_io_in_bits_Decode_cf_intrVec_11),
    .io_in_bits_Decode_cf_crossPageIPFFix(stage1_io_in_bits_Decode_cf_crossPageIPFFix),
    .io_in_bits_Decode_cf_runahead_checkpoint_id(stage1_io_in_bits_Decode_cf_runahead_checkpoint_id),
    .io_in_bits_Decode_ctrl_rfWen(stage1_io_in_bits_Decode_ctrl_rfWen),
    .io_in_bits_Decode_ctrl_rfDest(stage1_io_in_bits_Decode_ctrl_rfDest),
    .io_in_bits_Decode_ctrl_isMou(stage1_io_in_bits_Decode_ctrl_isMou),
    .io_in_bits_Decode_InstNo(stage1_io_in_bits_Decode_InstNo),
    .io_in_bits_Decode_InstFlag(stage1_io_in_bits_Decode_InstFlag),
    .io_in_bits_wdata(stage1_io_in_bits_wdata),
    .io_in_bits_src1(stage1_io_in_bits_src1),
    .io_in_bits_src2(stage1_io_in_bits_src2),
    .io_in_bits_func(stage1_io_in_bits_func),
    .io_out_ready(stage1_io_out_ready),
    .io_out_valid(stage1_io_out_valid),
    .io_out_bits_isMMIO(stage1_io_out_bits_isMMIO),
    .io_out_bits_loadAddrMisaligned(stage1_io_out_bits_loadAddrMisaligned),
    .io_out_bits_storeAddrMisaligned(stage1_io_out_bits_storeAddrMisaligned),
    .io_out_bits_Decode_cf_pc(stage1_io_out_bits_Decode_cf_pc),
    .io_out_bits_Decode_cf_exceptionVec_1(stage1_io_out_bits_Decode_cf_exceptionVec_1),
    .io_out_bits_Decode_cf_exceptionVec_2(stage1_io_out_bits_Decode_cf_exceptionVec_2),
    .io_out_bits_Decode_cf_exceptionVec_12(stage1_io_out_bits_Decode_cf_exceptionVec_12),
    .io_out_bits_Decode_cf_intrVec_0(stage1_io_out_bits_Decode_cf_intrVec_0),
    .io_out_bits_Decode_cf_intrVec_1(stage1_io_out_bits_Decode_cf_intrVec_1),
    .io_out_bits_Decode_cf_intrVec_2(stage1_io_out_bits_Decode_cf_intrVec_2),
    .io_out_bits_Decode_cf_intrVec_3(stage1_io_out_bits_Decode_cf_intrVec_3),
    .io_out_bits_Decode_cf_intrVec_4(stage1_io_out_bits_Decode_cf_intrVec_4),
    .io_out_bits_Decode_cf_intrVec_5(stage1_io_out_bits_Decode_cf_intrVec_5),
    .io_out_bits_Decode_cf_intrVec_6(stage1_io_out_bits_Decode_cf_intrVec_6),
    .io_out_bits_Decode_cf_intrVec_7(stage1_io_out_bits_Decode_cf_intrVec_7),
    .io_out_bits_Decode_cf_intrVec_8(stage1_io_out_bits_Decode_cf_intrVec_8),
    .io_out_bits_Decode_cf_intrVec_9(stage1_io_out_bits_Decode_cf_intrVec_9),
    .io_out_bits_Decode_cf_intrVec_10(stage1_io_out_bits_Decode_cf_intrVec_10),
    .io_out_bits_Decode_cf_intrVec_11(stage1_io_out_bits_Decode_cf_intrVec_11),
    .io_out_bits_Decode_cf_crossPageIPFFix(stage1_io_out_bits_Decode_cf_crossPageIPFFix),
    .io_out_bits_Decode_cf_runahead_checkpoint_id(stage1_io_out_bits_Decode_cf_runahead_checkpoint_id),
    .io_out_bits_Decode_ctrl_rfWen(stage1_io_out_bits_Decode_ctrl_rfWen),
    .io_out_bits_Decode_ctrl_rfDest(stage1_io_out_bits_Decode_ctrl_rfDest),
    .io_out_bits_Decode_ctrl_isMou(stage1_io_out_bits_Decode_ctrl_isMou),
    .io_out_bits_Decode_InstNo(stage1_io_out_bits_Decode_InstNo),
    .io_out_bits_Decode_InstFlag(stage1_io_out_bits_Decode_InstFlag),
    .io_out_bits_loadPF(stage1_io_out_bits_loadPF),
    .io_out_bits_storePF(stage1_io_out_bits_storePF),
    .io_out_bits_func(stage1_io_out_bits_func),
    .io_out_bits_addr(stage1_io_out_bits_addr),
    .io_dmem_req_ready(stage1_io_dmem_req_ready),
    .io_dmem_req_valid(stage1_io_dmem_req_valid),
    .io_dmem_req_bits_addr(stage1_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(stage1_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(stage1_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(stage1_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(stage1_io_dmem_req_bits_wdata),
    .io_flush(stage1_io_flush),
    .DTLBPF(stage1_DTLBPF),
    .loadPF_0(stage1_loadPF_0),
    .lsuMMIO_0(stage1_lsuMMIO_0),
    .storePF_0(stage1_storePF_0),
    .DTLBENABLE(stage1_DTLBENABLE),
    .DTLBFINISH(stage1_DTLBFINISH)
  );
  pipeline_lsu_stage2 stage2 ( // @[SIMD_PipeLSU.scala 653:22]
    .clock(stage2_clock),
    .reset(stage2_reset),
    .io_in_ready(stage2_io_in_ready),
    .io_in_valid(stage2_io_in_valid),
    .io_in_bits_isMMIO(stage2_io_in_bits_isMMIO),
    .io_in_bits_loadAddrMisaligned(stage2_io_in_bits_loadAddrMisaligned),
    .io_in_bits_storeAddrMisaligned(stage2_io_in_bits_storeAddrMisaligned),
    .io_in_bits_Decode_cf_pc(stage2_io_in_bits_Decode_cf_pc),
    .io_in_bits_Decode_cf_exceptionVec_1(stage2_io_in_bits_Decode_cf_exceptionVec_1),
    .io_in_bits_Decode_cf_exceptionVec_2(stage2_io_in_bits_Decode_cf_exceptionVec_2),
    .io_in_bits_Decode_cf_exceptionVec_12(stage2_io_in_bits_Decode_cf_exceptionVec_12),
    .io_in_bits_Decode_cf_intrVec_0(stage2_io_in_bits_Decode_cf_intrVec_0),
    .io_in_bits_Decode_cf_intrVec_1(stage2_io_in_bits_Decode_cf_intrVec_1),
    .io_in_bits_Decode_cf_intrVec_2(stage2_io_in_bits_Decode_cf_intrVec_2),
    .io_in_bits_Decode_cf_intrVec_3(stage2_io_in_bits_Decode_cf_intrVec_3),
    .io_in_bits_Decode_cf_intrVec_4(stage2_io_in_bits_Decode_cf_intrVec_4),
    .io_in_bits_Decode_cf_intrVec_5(stage2_io_in_bits_Decode_cf_intrVec_5),
    .io_in_bits_Decode_cf_intrVec_6(stage2_io_in_bits_Decode_cf_intrVec_6),
    .io_in_bits_Decode_cf_intrVec_7(stage2_io_in_bits_Decode_cf_intrVec_7),
    .io_in_bits_Decode_cf_intrVec_8(stage2_io_in_bits_Decode_cf_intrVec_8),
    .io_in_bits_Decode_cf_intrVec_9(stage2_io_in_bits_Decode_cf_intrVec_9),
    .io_in_bits_Decode_cf_intrVec_10(stage2_io_in_bits_Decode_cf_intrVec_10),
    .io_in_bits_Decode_cf_intrVec_11(stage2_io_in_bits_Decode_cf_intrVec_11),
    .io_in_bits_Decode_cf_crossPageIPFFix(stage2_io_in_bits_Decode_cf_crossPageIPFFix),
    .io_in_bits_Decode_cf_runahead_checkpoint_id(stage2_io_in_bits_Decode_cf_runahead_checkpoint_id),
    .io_in_bits_Decode_ctrl_rfWen(stage2_io_in_bits_Decode_ctrl_rfWen),
    .io_in_bits_Decode_ctrl_rfDest(stage2_io_in_bits_Decode_ctrl_rfDest),
    .io_in_bits_Decode_ctrl_isMou(stage2_io_in_bits_Decode_ctrl_isMou),
    .io_in_bits_Decode_InstNo(stage2_io_in_bits_Decode_InstNo),
    .io_in_bits_Decode_InstFlag(stage2_io_in_bits_Decode_InstFlag),
    .io_in_bits_loadPF(stage2_io_in_bits_loadPF),
    .io_in_bits_storePF(stage2_io_in_bits_storePF),
    .io_in_bits_func(stage2_io_in_bits_func),
    .io_in_bits_addr(stage2_io_in_bits_addr),
    .io_out_ready(stage2_io_out_ready),
    .io_out_valid(stage2_io_out_valid),
    .io_out_bits_isMMIO(stage2_io_out_bits_isMMIO),
    .io_out_bits_loadAddrMisaligned(stage2_io_out_bits_loadAddrMisaligned),
    .io_out_bits_storeAddrMisaligned(stage2_io_out_bits_storeAddrMisaligned),
    .io_out_bits_Decode_cf_pc(stage2_io_out_bits_Decode_cf_pc),
    .io_out_bits_Decode_cf_exceptionVec_1(stage2_io_out_bits_Decode_cf_exceptionVec_1),
    .io_out_bits_Decode_cf_exceptionVec_2(stage2_io_out_bits_Decode_cf_exceptionVec_2),
    .io_out_bits_Decode_cf_exceptionVec_12(stage2_io_out_bits_Decode_cf_exceptionVec_12),
    .io_out_bits_Decode_cf_intrVec_0(stage2_io_out_bits_Decode_cf_intrVec_0),
    .io_out_bits_Decode_cf_intrVec_1(stage2_io_out_bits_Decode_cf_intrVec_1),
    .io_out_bits_Decode_cf_intrVec_2(stage2_io_out_bits_Decode_cf_intrVec_2),
    .io_out_bits_Decode_cf_intrVec_3(stage2_io_out_bits_Decode_cf_intrVec_3),
    .io_out_bits_Decode_cf_intrVec_4(stage2_io_out_bits_Decode_cf_intrVec_4),
    .io_out_bits_Decode_cf_intrVec_5(stage2_io_out_bits_Decode_cf_intrVec_5),
    .io_out_bits_Decode_cf_intrVec_6(stage2_io_out_bits_Decode_cf_intrVec_6),
    .io_out_bits_Decode_cf_intrVec_7(stage2_io_out_bits_Decode_cf_intrVec_7),
    .io_out_bits_Decode_cf_intrVec_8(stage2_io_out_bits_Decode_cf_intrVec_8),
    .io_out_bits_Decode_cf_intrVec_9(stage2_io_out_bits_Decode_cf_intrVec_9),
    .io_out_bits_Decode_cf_intrVec_10(stage2_io_out_bits_Decode_cf_intrVec_10),
    .io_out_bits_Decode_cf_intrVec_11(stage2_io_out_bits_Decode_cf_intrVec_11),
    .io_out_bits_Decode_cf_crossPageIPFFix(stage2_io_out_bits_Decode_cf_crossPageIPFFix),
    .io_out_bits_Decode_cf_runahead_checkpoint_id(stage2_io_out_bits_Decode_cf_runahead_checkpoint_id),
    .io_out_bits_Decode_ctrl_rfWen(stage2_io_out_bits_Decode_ctrl_rfWen),
    .io_out_bits_Decode_ctrl_rfDest(stage2_io_out_bits_Decode_ctrl_rfDest),
    .io_out_bits_Decode_ctrl_isMou(stage2_io_out_bits_Decode_ctrl_isMou),
    .io_out_bits_Decode_InstNo(stage2_io_out_bits_Decode_InstNo),
    .io_out_bits_Decode_InstFlag(stage2_io_out_bits_Decode_InstFlag),
    .io_out_bits_loadPF(stage2_io_out_bits_loadPF),
    .io_out_bits_storePF(stage2_io_out_bits_storePF),
    .io_out_bits_result(stage2_io_out_bits_result),
    .io_out_bits_addr(stage2_io_out_bits_addr),
    .io_dmem_req_valid(stage2_io_dmem_req_valid),
    .io_dmem_req_bits_cmd(stage2_io_dmem_req_bits_cmd),
    .io_dmem_resp_ready(stage2_io_dmem_resp_ready),
    .io_dmem_resp_valid(stage2_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(stage2_io_dmem_resp_bits_rdata),
    .io_flush(stage2_io_flush)
  );
  pipeline_lsu_empty_stage stage_empty ( // @[SIMD_PipeLSU.scala 654:27]
    .io_in_ready(stage_empty_io_in_ready),
    .io_in_valid(stage_empty_io_in_valid),
    .io_in_bits_loadAddrMisaligned(stage_empty_io_in_bits_loadAddrMisaligned),
    .io_in_bits_storeAddrMisaligned(stage_empty_io_in_bits_storeAddrMisaligned),
    .io_in_bits_Decode_cf_pc(stage_empty_io_in_bits_Decode_cf_pc),
    .io_in_bits_Decode_cf_exceptionVec_1(stage_empty_io_in_bits_Decode_cf_exceptionVec_1),
    .io_in_bits_Decode_cf_exceptionVec_2(stage_empty_io_in_bits_Decode_cf_exceptionVec_2),
    .io_in_bits_Decode_cf_exceptionVec_12(stage_empty_io_in_bits_Decode_cf_exceptionVec_12),
    .io_in_bits_Decode_cf_intrVec_0(stage_empty_io_in_bits_Decode_cf_intrVec_0),
    .io_in_bits_Decode_cf_intrVec_1(stage_empty_io_in_bits_Decode_cf_intrVec_1),
    .io_in_bits_Decode_cf_intrVec_2(stage_empty_io_in_bits_Decode_cf_intrVec_2),
    .io_in_bits_Decode_cf_intrVec_3(stage_empty_io_in_bits_Decode_cf_intrVec_3),
    .io_in_bits_Decode_cf_intrVec_4(stage_empty_io_in_bits_Decode_cf_intrVec_4),
    .io_in_bits_Decode_cf_intrVec_5(stage_empty_io_in_bits_Decode_cf_intrVec_5),
    .io_in_bits_Decode_cf_intrVec_6(stage_empty_io_in_bits_Decode_cf_intrVec_6),
    .io_in_bits_Decode_cf_intrVec_7(stage_empty_io_in_bits_Decode_cf_intrVec_7),
    .io_in_bits_Decode_cf_intrVec_8(stage_empty_io_in_bits_Decode_cf_intrVec_8),
    .io_in_bits_Decode_cf_intrVec_9(stage_empty_io_in_bits_Decode_cf_intrVec_9),
    .io_in_bits_Decode_cf_intrVec_10(stage_empty_io_in_bits_Decode_cf_intrVec_10),
    .io_in_bits_Decode_cf_intrVec_11(stage_empty_io_in_bits_Decode_cf_intrVec_11),
    .io_in_bits_Decode_cf_crossPageIPFFix(stage_empty_io_in_bits_Decode_cf_crossPageIPFFix),
    .io_in_bits_Decode_cf_runahead_checkpoint_id(stage_empty_io_in_bits_Decode_cf_runahead_checkpoint_id),
    .io_in_bits_Decode_ctrl_rfWen(stage_empty_io_in_bits_Decode_ctrl_rfWen),
    .io_in_bits_Decode_ctrl_rfDest(stage_empty_io_in_bits_Decode_ctrl_rfDest),
    .io_in_bits_Decode_ctrl_isMou(stage_empty_io_in_bits_Decode_ctrl_isMou),
    .io_in_bits_Decode_InstNo(stage_empty_io_in_bits_Decode_InstNo),
    .io_in_bits_Decode_InstFlag(stage_empty_io_in_bits_Decode_InstFlag),
    .io_in_bits_loadPF(stage_empty_io_in_bits_loadPF),
    .io_in_bits_storePF(stage_empty_io_in_bits_storePF),
    .io_in_bits_result(stage_empty_io_in_bits_result),
    .io_in_bits_addr(stage_empty_io_in_bits_addr),
    .io_out_ready(stage_empty_io_out_ready),
    .io_out_valid(stage_empty_io_out_valid),
    .io_out_bits_loadAddrMisaligned(stage_empty_io_out_bits_loadAddrMisaligned),
    .io_out_bits_storeAddrMisaligned(stage_empty_io_out_bits_storeAddrMisaligned),
    .io_out_bits_Decode_cf_pc(stage_empty_io_out_bits_Decode_cf_pc),
    .io_out_bits_Decode_cf_exceptionVec_1(stage_empty_io_out_bits_Decode_cf_exceptionVec_1),
    .io_out_bits_Decode_cf_exceptionVec_2(stage_empty_io_out_bits_Decode_cf_exceptionVec_2),
    .io_out_bits_Decode_cf_exceptionVec_12(stage_empty_io_out_bits_Decode_cf_exceptionVec_12),
    .io_out_bits_Decode_cf_intrVec_0(stage_empty_io_out_bits_Decode_cf_intrVec_0),
    .io_out_bits_Decode_cf_intrVec_1(stage_empty_io_out_bits_Decode_cf_intrVec_1),
    .io_out_bits_Decode_cf_intrVec_2(stage_empty_io_out_bits_Decode_cf_intrVec_2),
    .io_out_bits_Decode_cf_intrVec_3(stage_empty_io_out_bits_Decode_cf_intrVec_3),
    .io_out_bits_Decode_cf_intrVec_4(stage_empty_io_out_bits_Decode_cf_intrVec_4),
    .io_out_bits_Decode_cf_intrVec_5(stage_empty_io_out_bits_Decode_cf_intrVec_5),
    .io_out_bits_Decode_cf_intrVec_6(stage_empty_io_out_bits_Decode_cf_intrVec_6),
    .io_out_bits_Decode_cf_intrVec_7(stage_empty_io_out_bits_Decode_cf_intrVec_7),
    .io_out_bits_Decode_cf_intrVec_8(stage_empty_io_out_bits_Decode_cf_intrVec_8),
    .io_out_bits_Decode_cf_intrVec_9(stage_empty_io_out_bits_Decode_cf_intrVec_9),
    .io_out_bits_Decode_cf_intrVec_10(stage_empty_io_out_bits_Decode_cf_intrVec_10),
    .io_out_bits_Decode_cf_intrVec_11(stage_empty_io_out_bits_Decode_cf_intrVec_11),
    .io_out_bits_Decode_cf_crossPageIPFFix(stage_empty_io_out_bits_Decode_cf_crossPageIPFFix),
    .io_out_bits_Decode_cf_runahead_checkpoint_id(stage_empty_io_out_bits_Decode_cf_runahead_checkpoint_id),
    .io_out_bits_Decode_ctrl_rfWen(stage_empty_io_out_bits_Decode_ctrl_rfWen),
    .io_out_bits_Decode_ctrl_rfDest(stage_empty_io_out_bits_Decode_ctrl_rfDest),
    .io_out_bits_Decode_ctrl_isMou(stage_empty_io_out_bits_Decode_ctrl_isMou),
    .io_out_bits_Decode_InstNo(stage_empty_io_out_bits_Decode_InstNo),
    .io_out_bits_Decode_InstFlag(stage_empty_io_out_bits_Decode_InstFlag),
    .io_out_bits_loadPF(stage_empty_io_out_bits_loadPF),
    .io_out_bits_storePF(stage_empty_io_out_bits_storePF),
    .io_out_bits_result(stage_empty_io_out_bits_result),
    .io_out_bits_addr(stage_empty_io_out_bits_addr)
  );
  lsu_for_atom atomstage ( // @[SIMD_PipeLSU.scala 655:25]
    .clock(atomstage_clock),
    .reset(atomstage_reset),
    .io_in_valid(atomstage_io_in_valid),
    .io_in_bits_Decode_cf_instr(atomstage_io_in_bits_Decode_cf_instr),
    .io_in_bits_Decode_cf_pc(atomstage_io_in_bits_Decode_cf_pc),
    .io_in_bits_Decode_cf_exceptionVec_1(atomstage_io_in_bits_Decode_cf_exceptionVec_1),
    .io_in_bits_Decode_cf_exceptionVec_2(atomstage_io_in_bits_Decode_cf_exceptionVec_2),
    .io_in_bits_Decode_cf_exceptionVec_12(atomstage_io_in_bits_Decode_cf_exceptionVec_12),
    .io_in_bits_Decode_cf_intrVec_0(atomstage_io_in_bits_Decode_cf_intrVec_0),
    .io_in_bits_Decode_cf_intrVec_1(atomstage_io_in_bits_Decode_cf_intrVec_1),
    .io_in_bits_Decode_cf_intrVec_2(atomstage_io_in_bits_Decode_cf_intrVec_2),
    .io_in_bits_Decode_cf_intrVec_3(atomstage_io_in_bits_Decode_cf_intrVec_3),
    .io_in_bits_Decode_cf_intrVec_4(atomstage_io_in_bits_Decode_cf_intrVec_4),
    .io_in_bits_Decode_cf_intrVec_5(atomstage_io_in_bits_Decode_cf_intrVec_5),
    .io_in_bits_Decode_cf_intrVec_6(atomstage_io_in_bits_Decode_cf_intrVec_6),
    .io_in_bits_Decode_cf_intrVec_7(atomstage_io_in_bits_Decode_cf_intrVec_7),
    .io_in_bits_Decode_cf_intrVec_8(atomstage_io_in_bits_Decode_cf_intrVec_8),
    .io_in_bits_Decode_cf_intrVec_9(atomstage_io_in_bits_Decode_cf_intrVec_9),
    .io_in_bits_Decode_cf_intrVec_10(atomstage_io_in_bits_Decode_cf_intrVec_10),
    .io_in_bits_Decode_cf_intrVec_11(atomstage_io_in_bits_Decode_cf_intrVec_11),
    .io_in_bits_Decode_cf_crossPageIPFFix(atomstage_io_in_bits_Decode_cf_crossPageIPFFix),
    .io_in_bits_Decode_cf_runahead_checkpoint_id(atomstage_io_in_bits_Decode_cf_runahead_checkpoint_id),
    .io_in_bits_Decode_ctrl_rfWen(atomstage_io_in_bits_Decode_ctrl_rfWen),
    .io_in_bits_Decode_ctrl_rfDest(atomstage_io_in_bits_Decode_ctrl_rfDest),
    .io_in_bits_Decode_ctrl_isMou(atomstage_io_in_bits_Decode_ctrl_isMou),
    .io_in_bits_Decode_InstNo(atomstage_io_in_bits_Decode_InstNo),
    .io_in_bits_Decode_InstFlag(atomstage_io_in_bits_Decode_InstFlag),
    .io_in_bits_wdata(atomstage_io_in_bits_wdata),
    .io_in_bits_src1(atomstage_io_in_bits_src1),
    .io_in_bits_src2(atomstage_io_in_bits_src2),
    .io_in_bits_func(atomstage_io_in_bits_func),
    .io_out_ready(atomstage_io_out_ready),
    .io_out_valid(atomstage_io_out_valid),
    .io_out_bits_loadAddrMisaligned(atomstage_io_out_bits_loadAddrMisaligned),
    .io_out_bits_storeAddrMisaligned(atomstage_io_out_bits_storeAddrMisaligned),
    .io_out_bits_Decode_cf_pc(atomstage_io_out_bits_Decode_cf_pc),
    .io_out_bits_Decode_cf_exceptionVec_1(atomstage_io_out_bits_Decode_cf_exceptionVec_1),
    .io_out_bits_Decode_cf_exceptionVec_2(atomstage_io_out_bits_Decode_cf_exceptionVec_2),
    .io_out_bits_Decode_cf_exceptionVec_12(atomstage_io_out_bits_Decode_cf_exceptionVec_12),
    .io_out_bits_Decode_cf_intrVec_0(atomstage_io_out_bits_Decode_cf_intrVec_0),
    .io_out_bits_Decode_cf_intrVec_1(atomstage_io_out_bits_Decode_cf_intrVec_1),
    .io_out_bits_Decode_cf_intrVec_2(atomstage_io_out_bits_Decode_cf_intrVec_2),
    .io_out_bits_Decode_cf_intrVec_3(atomstage_io_out_bits_Decode_cf_intrVec_3),
    .io_out_bits_Decode_cf_intrVec_4(atomstage_io_out_bits_Decode_cf_intrVec_4),
    .io_out_bits_Decode_cf_intrVec_5(atomstage_io_out_bits_Decode_cf_intrVec_5),
    .io_out_bits_Decode_cf_intrVec_6(atomstage_io_out_bits_Decode_cf_intrVec_6),
    .io_out_bits_Decode_cf_intrVec_7(atomstage_io_out_bits_Decode_cf_intrVec_7),
    .io_out_bits_Decode_cf_intrVec_8(atomstage_io_out_bits_Decode_cf_intrVec_8),
    .io_out_bits_Decode_cf_intrVec_9(atomstage_io_out_bits_Decode_cf_intrVec_9),
    .io_out_bits_Decode_cf_intrVec_10(atomstage_io_out_bits_Decode_cf_intrVec_10),
    .io_out_bits_Decode_cf_intrVec_11(atomstage_io_out_bits_Decode_cf_intrVec_11),
    .io_out_bits_Decode_cf_crossPageIPFFix(atomstage_io_out_bits_Decode_cf_crossPageIPFFix),
    .io_out_bits_Decode_cf_runahead_checkpoint_id(atomstage_io_out_bits_Decode_cf_runahead_checkpoint_id),
    .io_out_bits_Decode_ctrl_rfWen(atomstage_io_out_bits_Decode_ctrl_rfWen),
    .io_out_bits_Decode_ctrl_rfDest(atomstage_io_out_bits_Decode_ctrl_rfDest),
    .io_out_bits_Decode_ctrl_isMou(atomstage_io_out_bits_Decode_ctrl_isMou),
    .io_out_bits_Decode_InstNo(atomstage_io_out_bits_Decode_InstNo),
    .io_out_bits_Decode_InstFlag(atomstage_io_out_bits_Decode_InstFlag),
    .io_out_bits_loadPF(atomstage_io_out_bits_loadPF),
    .io_out_bits_storePF(atomstage_io_out_bits_storePF),
    .io_out_bits_result(atomstage_io_out_bits_result),
    .io_dmem_req_ready(atomstage_io_dmem_req_ready),
    .io_dmem_req_valid(atomstage_io_dmem_req_valid),
    .io_dmem_req_bits_addr(atomstage_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(atomstage_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(atomstage_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(atomstage_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(atomstage_io_dmem_req_bits_wdata),
    .io_dmem_resp_ready(atomstage_io_dmem_resp_ready),
    .io_dmem_resp_valid(atomstage_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(atomstage_io_dmem_resp_bits_rdata),
    .io_flush(atomstage_io_flush),
    .setLr_0(atomstage_setLr_0),
    .DTLBPF(atomstage_DTLBPF),
    .loadPF_0(atomstage_loadPF_0),
    .lr_0(atomstage_lr_0),
    .amoReq_0(atomstage_amoReq_0),
    .storePF_0(atomstage_storePF_0),
    .DTLBENABLE(atomstage_DTLBENABLE),
    .DTLBFINISH(atomstage_DTLBFINISH),
    .setLrAddr_0(atomstage_setLrAddr_0),
    .setLrVal_0(atomstage_setLrVal_0),
    .lr_addr(atomstage_lr_addr)
  );
  assign io_in_ready = ~io_in_valid | lsu_firststage_fire; // @[SIMD_PipeLSU.scala 742:26]
  assign io_out_valid = stage_empty_io_in_valid ? stage_empty_io_out_valid : stage2_io_out_valid & _T; // @[SIMD_PipeLSU.scala 719:32 720:17 725:17]
  assign io_out_bits = stage_empty_io_in_valid ? stage_empty_io_out_bits_result : stage2_io_out_bits_result; // @[SIMD_PipeLSU.scala 719:32 721:17 726:17]
  assign io_dmem_req_valid = atomstage_io_in_valid ? atomstage_io_dmem_req_valid : stage1_io_dmem_req_valid; // @[SIMD_PipeLSU.scala 731:30 732:13 735:17]
  assign io_dmem_req_bits_addr = atomstage_io_in_valid ? atomstage_io_dmem_req_bits_addr : stage1_io_dmem_req_bits_addr; // @[SIMD_PipeLSU.scala 731:30 732:13 735:17]
  assign io_dmem_req_bits_size = atomstage_io_in_valid ? atomstage_io_dmem_req_bits_size : stage1_io_dmem_req_bits_size; // @[SIMD_PipeLSU.scala 731:30 732:13 735:17]
  assign io_dmem_req_bits_cmd = atomstage_io_in_valid ? atomstage_io_dmem_req_bits_cmd : stage1_io_dmem_req_bits_cmd; // @[SIMD_PipeLSU.scala 731:30 732:13 735:17]
  assign io_dmem_req_bits_wmask = atomstage_io_in_valid ? atomstage_io_dmem_req_bits_wmask :
    stage1_io_dmem_req_bits_wmask; // @[SIMD_PipeLSU.scala 731:30 732:13 735:17]
  assign io_dmem_req_bits_wdata = atomstage_io_in_valid ? atomstage_io_dmem_req_bits_wdata :
    stage1_io_dmem_req_bits_wdata; // @[SIMD_PipeLSU.scala 731:30 732:13 735:17]
  assign io_loadAddrMisaligned = stage_empty_io_out_valid & stage_empty_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 714:54]
  assign io_storeAddrMisaligned = stage_empty_io_out_valid & stage_empty_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 715:54]
  assign io_DecodeOut_cf_pc = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_pc :
    stage2_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_exceptionVec_1 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_exceptionVec_1 :
    stage2_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_exceptionVec_2 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_exceptionVec_2 :
    stage2_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_exceptionVec_12 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_exceptionVec_12
     : stage2_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_0 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_0 :
    stage2_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_1 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_1 :
    stage2_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_2 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_2 :
    stage2_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_3 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_3 :
    stage2_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_4 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_4 :
    stage2_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_5 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_5 :
    stage2_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_6 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_6 :
    stage2_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_7 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_7 :
    stage2_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_8 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_8 :
    stage2_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_9 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_9 :
    stage2_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_10 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_10 :
    stage2_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_intrVec_11 = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_intrVec_11 :
    stage2_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_crossPageIPFFix = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_cf_crossPageIPFFix
     : stage2_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_cf_runahead_checkpoint_id = stage_empty_io_in_valid ?
    stage_empty_io_out_bits_Decode_cf_runahead_checkpoint_id : stage2_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_ctrl_rfWen = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_ctrl_rfWen :
    stage2_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_ctrl_rfDest = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_ctrl_rfDest :
    stage2_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_ctrl_isMou = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_ctrl_isMou :
    stage2_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_InstNo = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_InstNo :
    stage2_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_DecodeOut_InstFlag = stage_empty_io_in_valid ? stage_empty_io_out_bits_Decode_InstFlag :
    stage2_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 719:32 723:17 728:17]
  assign io_loadPF = stage_empty_io_out_valid & stage_empty_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 717:43]
  assign io_storePF = stage_empty_io_out_valid & stage_empty_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 716:43]
  assign lsu_firststage_fire_0 = lsu_firststage_fire;
  assign setLr = atomstage_setLr_0;
  assign amoReq = atomstage_amoReq_0;
  assign addr_0 = addr;
  assign setLrAddr = atomstage_setLrAddr_0;
  assign setLrVal = atomstage_setLrVal_0;
  assign stage1_clock = clock;
  assign stage1_reset = reset;
  assign stage1_io_in_valid = io_in_valid & ~stage2_exp & ~stage_empty_exp & ~atomReq & _T_6; // @[SIMD_PipeLSU.scala 667:78]
  assign stage1_io_in_bits_Decode_cf_pc = io_DecodeIn_cf_pc; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_exceptionVec_1 = io_DecodeIn_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_exceptionVec_2 = io_DecodeIn_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_exceptionVec_12 = io_DecodeIn_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_0 = io_DecodeIn_cf_intrVec_0; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_1 = io_DecodeIn_cf_intrVec_1; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_2 = io_DecodeIn_cf_intrVec_2; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_3 = io_DecodeIn_cf_intrVec_3; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_4 = io_DecodeIn_cf_intrVec_4; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_5 = io_DecodeIn_cf_intrVec_5; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_6 = io_DecodeIn_cf_intrVec_6; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_7 = io_DecodeIn_cf_intrVec_7; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_8 = io_DecodeIn_cf_intrVec_8; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_9 = io_DecodeIn_cf_intrVec_9; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_10 = io_DecodeIn_cf_intrVec_10; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_intrVec_11 = io_DecodeIn_cf_intrVec_11; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_crossPageIPFFix = io_DecodeIn_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_cf_runahead_checkpoint_id = io_DecodeIn_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_ctrl_rfWen = io_DecodeIn_ctrl_rfWen; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_ctrl_rfDest = io_DecodeIn_ctrl_rfDest; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_ctrl_isMou = io_DecodeIn_ctrl_isMou; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_InstNo = io_DecodeIn_InstNo; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_Decode_InstFlag = io_DecodeIn_InstFlag; // @[SIMD_PipeLSU.scala 674:27]
  assign stage1_io_in_bits_wdata = io_wdata; // @[SIMD_PipeLSU.scala 673:27]
  assign stage1_io_in_bits_src1 = io_in_bits_src1; // @[SIMD_PipeLSU.scala 670:27]
  assign stage1_io_in_bits_src2 = io_in_bits_src2; // @[SIMD_PipeLSU.scala 671:27]
  assign stage1_io_in_bits_func = io_in_bits_func; // @[SIMD_PipeLSU.scala 672:27]
  assign stage1_io_out_ready = stage2_io_in_ready; // @[Pipeline.scala 29:16]
  assign stage1_io_dmem_req_ready = atomstage_io_in_valid ? 1'h0 : io_dmem_req_ready; // @[SIMD_PipeLSU.scala 698:18 731:30 735:17]
  assign stage1_io_flush = io_flush; // @[SIMD_PipeLSU.scala 668:22]
  assign stage1_DTLBPF = _T_408;
  assign stage1_loadPF_0 = io_memMMU_dmem_loadPF;
  assign stage1_lsuMMIO_0 = ismmio;
  assign stage1_storePF_0 = io_memMMU_dmem_storePF;
  assign stage1_DTLBENABLE = vmEnable;
  assign stage1_DTLBFINISH = _T_407;
  assign stage2_clock = clock;
  assign stage2_reset = reset;
  assign stage2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign stage2_io_in_bits_isMMIO = r_isMMIO; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_loadAddrMisaligned = r_loadAddrMisaligned; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_storeAddrMisaligned = r_storeAddrMisaligned; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_pc = r_Decode_cf_pc; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_exceptionVec_1 = r_Decode_cf_exceptionVec_1; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_exceptionVec_2 = r_Decode_cf_exceptionVec_2; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_exceptionVec_12 = r_Decode_cf_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_0 = r_Decode_cf_intrVec_0; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_1 = r_Decode_cf_intrVec_1; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_2 = r_Decode_cf_intrVec_2; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_3 = r_Decode_cf_intrVec_3; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_4 = r_Decode_cf_intrVec_4; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_5 = r_Decode_cf_intrVec_5; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_6 = r_Decode_cf_intrVec_6; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_7 = r_Decode_cf_intrVec_7; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_8 = r_Decode_cf_intrVec_8; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_9 = r_Decode_cf_intrVec_9; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_10 = r_Decode_cf_intrVec_10; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_intrVec_11 = r_Decode_cf_intrVec_11; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_crossPageIPFFix = r_Decode_cf_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_cf_runahead_checkpoint_id = r_Decode_cf_runahead_checkpoint_id; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_ctrl_rfWen = r_Decode_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_ctrl_rfDest = r_Decode_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_ctrl_isMou = r_Decode_ctrl_isMou; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_InstNo = r_Decode_InstNo; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_Decode_InstFlag = r_Decode_InstFlag; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_loadPF = r_loadPF; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_storePF = r_storePF; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_func = r_func; // @[Pipeline.scala 30:16]
  assign stage2_io_in_bits_addr = r_addr; // @[Pipeline.scala 30:16]
  assign stage2_io_out_ready = atomstage_io_in_valid ? io_out_ready : _GEN_158; // @[SIMD_PipeLSU.scala 689:23 703:30]
  assign stage2_io_dmem_resp_valid = atomstage_io_in_valid ? 1'h0 : io_dmem_resp_valid; // @[SIMD_PipeLSU.scala 699:18 731:30 736:18]
  assign stage2_io_dmem_resp_bits_rdata = atomstage_io_in_valid ? 64'h0 : io_dmem_resp_bits_rdata; // @[SIMD_PipeLSU.scala 699:18 731:30 736:18]
  assign stage2_io_flush = io_flush; // @[SIMD_PipeLSU.scala 688:19]
  assign stage_empty_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign stage_empty_io_in_bits_loadAddrMisaligned = r_1_loadAddrMisaligned; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_storeAddrMisaligned = r_1_storeAddrMisaligned; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_pc = r_1_Decode_cf_pc; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_exceptionVec_1 = r_1_Decode_cf_exceptionVec_1; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_exceptionVec_2 = r_1_Decode_cf_exceptionVec_2; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_exceptionVec_12 = r_1_Decode_cf_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_0 = r_1_Decode_cf_intrVec_0; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_1 = r_1_Decode_cf_intrVec_1; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_2 = r_1_Decode_cf_intrVec_2; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_3 = r_1_Decode_cf_intrVec_3; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_4 = r_1_Decode_cf_intrVec_4; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_5 = r_1_Decode_cf_intrVec_5; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_6 = r_1_Decode_cf_intrVec_6; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_7 = r_1_Decode_cf_intrVec_7; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_8 = r_1_Decode_cf_intrVec_8; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_9 = r_1_Decode_cf_intrVec_9; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_10 = r_1_Decode_cf_intrVec_10; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_intrVec_11 = r_1_Decode_cf_intrVec_11; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_crossPageIPFFix = r_1_Decode_cf_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_cf_runahead_checkpoint_id = r_1_Decode_cf_runahead_checkpoint_id; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_ctrl_rfWen = r_1_Decode_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_ctrl_rfDest = r_1_Decode_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_ctrl_isMou = r_1_Decode_ctrl_isMou; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_InstNo = r_1_Decode_InstNo; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_Decode_InstFlag = r_1_Decode_InstFlag; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_loadPF = r_1_loadPF; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_storePF = r_1_storePF; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_result = r_1_result; // @[Pipeline.scala 30:16]
  assign stage_empty_io_in_bits_addr = r_1_addr; // @[Pipeline.scala 30:16]
  assign stage_empty_io_out_ready = io_out_ready; // @[SIMD_PipeLSU.scala 693:28]
  assign atomstage_clock = clock;
  assign atomstage_reset = reset;
  assign atomstage_io_in_valid = io_in_valid & atomReq & ~stage2_io_in_valid; // @[SIMD_PipeLSU.scala 676:45]
  assign atomstage_io_in_bits_Decode_cf_instr = io_DecodeIn_cf_instr; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_pc = io_DecodeIn_cf_pc; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_exceptionVec_1 = io_DecodeIn_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_exceptionVec_2 = io_DecodeIn_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_exceptionVec_12 = io_DecodeIn_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_0 = io_DecodeIn_cf_intrVec_0; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_1 = io_DecodeIn_cf_intrVec_1; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_2 = io_DecodeIn_cf_intrVec_2; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_3 = io_DecodeIn_cf_intrVec_3; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_4 = io_DecodeIn_cf_intrVec_4; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_5 = io_DecodeIn_cf_intrVec_5; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_6 = io_DecodeIn_cf_intrVec_6; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_7 = io_DecodeIn_cf_intrVec_7; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_8 = io_DecodeIn_cf_intrVec_8; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_9 = io_DecodeIn_cf_intrVec_9; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_10 = io_DecodeIn_cf_intrVec_10; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_intrVec_11 = io_DecodeIn_cf_intrVec_11; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_crossPageIPFFix = io_DecodeIn_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_cf_runahead_checkpoint_id = io_DecodeIn_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_ctrl_rfWen = io_DecodeIn_ctrl_rfWen; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_ctrl_rfDest = io_DecodeIn_ctrl_rfDest; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_ctrl_isMou = io_DecodeIn_ctrl_isMou; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_InstNo = io_DecodeIn_InstNo; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_Decode_InstFlag = io_DecodeIn_InstFlag; // @[SIMD_PipeLSU.scala 683:30]
  assign atomstage_io_in_bits_wdata = io_wdata; // @[SIMD_PipeLSU.scala 682:30]
  assign atomstage_io_in_bits_src1 = io_in_bits_src1; // @[SIMD_PipeLSU.scala 679:30]
  assign atomstage_io_in_bits_src2 = io_in_bits_src2; // @[SIMD_PipeLSU.scala 680:30]
  assign atomstage_io_in_bits_func = io_in_bits_func; // @[SIMD_PipeLSU.scala 681:30]
  assign atomstage_io_out_ready = atomstage_io_in_valid ? empty_out_ready : io_out_ready; // @[SIMD_PipeLSU.scala 703:30 706:28 684:30]
  assign atomstage_io_dmem_req_ready = atomstage_io_in_valid & io_dmem_req_ready; // @[SIMD_PipeLSU.scala 731:30 732:13 697:21]
  assign atomstage_io_dmem_resp_valid = atomstage_io_in_valid & io_dmem_resp_valid; // @[SIMD_PipeLSU.scala 731:30 732:13 697:21]
  assign atomstage_io_dmem_resp_bits_rdata = atomstage_io_in_valid ? io_dmem_resp_bits_rdata : 64'h0; // @[SIMD_PipeLSU.scala 731:30 732:13 697:21]
  assign atomstage_io_flush = io_flush; // @[SIMD_PipeLSU.scala 677:25]
  assign atomstage_DTLBPF = _T_408;
  assign atomstage_loadPF_0 = io_memMMU_dmem_loadPF;
  assign atomstage_lr_0 = lr;
  assign atomstage_storePF_0 = io_memMMU_dmem_storePF;
  assign atomstage_DTLBENABLE = vmEnable;
  assign atomstage_DTLBFINISH = _T_407;
  assign atomstage_lr_addr = lrAddr;
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_isMMIO <= stage1_io_out_bits_isMMIO; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_loadAddrMisaligned <= stage1_io_out_bits_loadAddrMisaligned; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_storeAddrMisaligned <= stage1_io_out_bits_storeAddrMisaligned; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_pc <= stage1_io_out_bits_Decode_cf_pc; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_exceptionVec_1 <= stage1_io_out_bits_Decode_cf_exceptionVec_1; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_exceptionVec_2 <= stage1_io_out_bits_Decode_cf_exceptionVec_2; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_exceptionVec_12 <= stage1_io_out_bits_Decode_cf_exceptionVec_12; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_0 <= stage1_io_out_bits_Decode_cf_intrVec_0; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_1 <= stage1_io_out_bits_Decode_cf_intrVec_1; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_2 <= stage1_io_out_bits_Decode_cf_intrVec_2; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_3 <= stage1_io_out_bits_Decode_cf_intrVec_3; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_4 <= stage1_io_out_bits_Decode_cf_intrVec_4; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_5 <= stage1_io_out_bits_Decode_cf_intrVec_5; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_6 <= stage1_io_out_bits_Decode_cf_intrVec_6; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_7 <= stage1_io_out_bits_Decode_cf_intrVec_7; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_8 <= stage1_io_out_bits_Decode_cf_intrVec_8; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_9 <= stage1_io_out_bits_Decode_cf_intrVec_9; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_10 <= stage1_io_out_bits_Decode_cf_intrVec_10; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_intrVec_11 <= stage1_io_out_bits_Decode_cf_intrVec_11; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_crossPageIPFFix <= stage1_io_out_bits_Decode_cf_crossPageIPFFix; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_cf_runahead_checkpoint_id <= stage1_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_ctrl_rfWen <= stage1_io_out_bits_Decode_ctrl_rfWen; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_ctrl_rfDest <= stage1_io_out_bits_Decode_ctrl_rfDest; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_ctrl_isMou <= stage1_io_out_bits_Decode_ctrl_isMou; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_InstNo <= stage1_io_out_bits_Decode_InstNo; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_Decode_InstFlag <= stage1_io_out_bits_Decode_InstFlag; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_loadPF <= stage1_io_out_bits_loadPF; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_storePF <= stage1_io_out_bits_storePF; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_func <= stage1_io_out_bits_func; // @[Reg.scala 16:23]
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      r_addr <= stage1_io_out_bits_addr; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush) begin // @[Pipeline.scala 27:20]
      REG_1 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_1 <= _GEN_240;
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_loadAddrMisaligned <= atomstage_io_out_bits_loadAddrMisaligned; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_loadAddrMisaligned <= _GEN_156;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_storeAddrMisaligned <= atomstage_io_out_bits_storeAddrMisaligned; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_storeAddrMisaligned <= _GEN_155;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_pc <= atomstage_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 705:21]
      end else if (stage2_io_in_valid & stage2_exp) begin // @[SIMD_PipeLSU.scala 707:47]
        r_1_Decode_cf_pc <= stage2_io_out_bits_Decode_cf_pc; // @[SIMD_PipeLSU.scala 709:21]
      end else begin
        r_1_Decode_cf_pc <= 39'h0;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_exceptionVec_1 <= atomstage_io_out_bits_Decode_cf_exceptionVec_1; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_exceptionVec_1 <= _GEN_134;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_exceptionVec_2 <= atomstage_io_out_bits_Decode_cf_exceptionVec_2; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_exceptionVec_2 <= _GEN_135;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_exceptionVec_12 <= atomstage_io_out_bits_Decode_cf_exceptionVec_12; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_exceptionVec_12 <= _GEN_145;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_0 <= atomstage_io_out_bits_Decode_cf_intrVec_0; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_0 <= _GEN_121;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_1 <= atomstage_io_out_bits_Decode_cf_intrVec_1; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_1 <= _GEN_122;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_2 <= atomstage_io_out_bits_Decode_cf_intrVec_2; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_2 <= _GEN_123;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_3 <= atomstage_io_out_bits_Decode_cf_intrVec_3; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_3 <= _GEN_124;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_4 <= atomstage_io_out_bits_Decode_cf_intrVec_4; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_4 <= _GEN_125;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_5 <= atomstage_io_out_bits_Decode_cf_intrVec_5; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_5 <= _GEN_126;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_6 <= atomstage_io_out_bits_Decode_cf_intrVec_6; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_6 <= _GEN_127;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_7 <= atomstage_io_out_bits_Decode_cf_intrVec_7; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_7 <= _GEN_128;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_8 <= atomstage_io_out_bits_Decode_cf_intrVec_8; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_8 <= _GEN_129;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_9 <= atomstage_io_out_bits_Decode_cf_intrVec_9; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_9 <= _GEN_130;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_10 <= atomstage_io_out_bits_Decode_cf_intrVec_10; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_10 <= _GEN_131;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_intrVec_11 <= atomstage_io_out_bits_Decode_cf_intrVec_11; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_intrVec_11 <= _GEN_132;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_crossPageIPFFix <= atomstage_io_out_bits_Decode_cf_crossPageIPFFix; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_cf_crossPageIPFFix <= _GEN_118;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_cf_runahead_checkpoint_id <= atomstage_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 705:21]
      end else if (stage2_io_in_valid & stage2_exp) begin // @[SIMD_PipeLSU.scala 707:47]
        r_1_Decode_cf_runahead_checkpoint_id <= stage2_io_out_bits_Decode_cf_runahead_checkpoint_id; // @[SIMD_PipeLSU.scala 709:21]
      end else begin
        r_1_Decode_cf_runahead_checkpoint_id <= 64'h0;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_ctrl_rfWen <= atomstage_io_out_bits_Decode_ctrl_rfWen; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_ctrl_rfWen <= _GEN_104;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_ctrl_rfDest <= atomstage_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 705:21]
      end else if (stage2_io_in_valid & stage2_exp) begin // @[SIMD_PipeLSU.scala 707:47]
        r_1_Decode_ctrl_rfDest <= stage2_io_out_bits_Decode_ctrl_rfDest; // @[SIMD_PipeLSU.scala 709:21]
      end else begin
        r_1_Decode_ctrl_rfDest <= 5'h0;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_ctrl_isMou <= atomstage_io_out_bits_Decode_ctrl_isMou; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_ctrl_isMou <= _GEN_96;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_InstNo <= atomstage_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 705:21]
      end else if (stage2_io_in_valid & stage2_exp) begin // @[SIMD_PipeLSU.scala 707:47]
        r_1_Decode_InstNo <= stage2_io_out_bits_Decode_InstNo; // @[SIMD_PipeLSU.scala 709:21]
      end else begin
        r_1_Decode_InstNo <= 5'h0;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_Decode_InstFlag <= atomstage_io_out_bits_Decode_InstFlag; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_Decode_InstFlag <= _GEN_89;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_loadPF <= atomstage_io_out_bits_loadPF; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_loadPF <= _GEN_88;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_storePF <= atomstage_io_out_bits_storePF; // @[SIMD_PipeLSU.scala 705:21]
      end else begin
        r_1_storePF <= _GEN_87;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_result <= atomstage_io_out_bits_result; // @[SIMD_PipeLSU.scala 705:21]
      end else if (stage2_io_in_valid & stage2_exp) begin // @[SIMD_PipeLSU.scala 707:47]
        r_1_result <= stage2_io_out_bits_result; // @[SIMD_PipeLSU.scala 709:21]
      end else begin
        r_1_result <= 64'h0;
      end
    end
    if (_T_24) begin // @[Reg.scala 16:19]
      if (atomstage_io_in_valid) begin // @[SIMD_PipeLSU.scala 703:30]
        r_1_addr <= 64'h0; // @[SIMD_PipeLSU.scala 705:21]
      end else if (stage2_io_in_valid & stage2_exp) begin // @[SIMD_PipeLSU.scala 707:47]
        r_1_addr <= stage2_io_out_bits_addr; // @[SIMD_PipeLSU.scala 709:21]
      end else begin
        r_1_addr <= 64'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_isMMIO = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_loadAddrMisaligned = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_storeAddrMisaligned = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  r_Decode_cf_pc = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  r_Decode_cf_exceptionVec_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_Decode_cf_exceptionVec_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_Decode_cf_exceptionVec_12 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_Decode_cf_intrVec_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_Decode_cf_intrVec_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_Decode_cf_intrVec_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_Decode_cf_intrVec_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_Decode_cf_intrVec_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_Decode_cf_intrVec_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_Decode_cf_intrVec_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_Decode_cf_intrVec_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_Decode_cf_intrVec_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_Decode_cf_intrVec_9 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_Decode_cf_intrVec_10 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_Decode_cf_intrVec_11 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_Decode_cf_crossPageIPFFix = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  r_Decode_cf_runahead_checkpoint_id = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  r_Decode_ctrl_rfWen = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_Decode_ctrl_rfDest = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  r_Decode_ctrl_isMou = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_Decode_InstNo = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  r_Decode_InstFlag = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_loadPF = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_storePF = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_func = _RAND_29[6:0];
  _RAND_30 = {2{`RANDOM}};
  r_addr = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  REG_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_1_loadAddrMisaligned = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_1_storeAddrMisaligned = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  r_1_Decode_cf_pc = _RAND_34[38:0];
  _RAND_35 = {1{`RANDOM}};
  r_1_Decode_cf_exceptionVec_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_1_Decode_cf_exceptionVec_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_1_Decode_cf_exceptionVec_12 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_2 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_3 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_4 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_5 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_6 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_7 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_8 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_9 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_10 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  r_1_Decode_cf_intrVec_11 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  r_1_Decode_cf_crossPageIPFFix = _RAND_50[0:0];
  _RAND_51 = {2{`RANDOM}};
  r_1_Decode_cf_runahead_checkpoint_id = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  r_1_Decode_ctrl_rfWen = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_1_Decode_ctrl_rfDest = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  r_1_Decode_ctrl_isMou = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  r_1_Decode_InstNo = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  r_1_Decode_InstFlag = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_1_loadPF = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  r_1_storePF = _RAND_58[0:0];
  _RAND_59 = {2{`RANDOM}};
  r_1_result = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  r_1_addr = _RAND_60[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module new_SIMD_CSR(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  output [63:0] io_out_bits,
  input  [38:0] io_cfIn_pc,
  input         io_cfIn_exceptionVec_1,
  input         io_cfIn_exceptionVec_2,
  input         io_cfIn_exceptionVec_4,
  input         io_cfIn_exceptionVec_6,
  input         io_cfIn_exceptionVec_12,
  input         io_cfIn_exceptionVec_13,
  input         io_cfIn_exceptionVec_15,
  input         io_cfIn_intrVec_0,
  input         io_cfIn_intrVec_1,
  input         io_cfIn_intrVec_2,
  input         io_cfIn_intrVec_3,
  input         io_cfIn_intrVec_4,
  input         io_cfIn_intrVec_5,
  input         io_cfIn_intrVec_6,
  input         io_cfIn_intrVec_7,
  input         io_cfIn_intrVec_8,
  input         io_cfIn_intrVec_9,
  input         io_cfIn_intrVec_10,
  input         io_cfIn_intrVec_11,
  input         io_cfIn_crossPageIPFFix,
  input         io_ctrlIn_isMou,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         io_instrValid,
  output [1:0]  io_imemMMU_priviledgeMode,
  output [1:0]  io_dmemMMU_priviledgeMode,
  output        io_dmemMMU_status_sum,
  output        io_dmemMMU_status_mxr,
  input         io_dmemMMU_loadPF,
  input         io_dmemMMU_storePF,
  input  [38:0] io_dmemMMU_addr,
  output        io_wenFix,
  input         set_lr,
  output        flushICache_0,
  output [63:0] satp_0,
  output        lr_0,
  input         OVWEN_0,
  input         mtip,
  input         meip,
  input  [63:0] LSUADDR,
  output [63:0] intrVec_0,
  input         msip,
  input  [63:0] set_lr_addr,
  output        flushTLB_0,
  input         set_lr_val,
  output [63:0] lrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  reg  lr; // @[SIMD_CSR.scala 560:19]
  reg [63:0] lrAddr; // @[SIMD_CSR.scala 561:23]
  reg [63:0] mtvec; // @[SIMD_CSR.scala 575:22]
  reg [63:0] mcounteren; // @[SIMD_CSR.scala 576:27]
  reg [63:0] mcause; // @[SIMD_CSR.scala 577:23]
  reg [63:0] mtval; // @[SIMD_CSR.scala 578:22]
  reg [63:0] mepc; // @[SIMD_CSR.scala 579:17]
  reg [63:0] mie; // @[SIMD_CSR.scala 581:20]
  reg [63:0] mipReg; // @[SIMD_CSR.scala 583:24]
  reg [63:0] mstatus; // @[SIMD_CSR.scala 598:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[SIMD_CSR.scala 599:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[SIMD_CSR.scala 599:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[SIMD_CSR.scala 599:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[SIMD_CSR.scala 599:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[SIMD_CSR.scala 599:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[SIMD_CSR.scala 599:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[SIMD_CSR.scala 599:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[SIMD_CSR.scala 599:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[SIMD_CSR.scala 599:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[SIMD_CSR.scala 599:39]
  reg [63:0] medeleg; // @[SIMD_CSR.scala 600:24]
  reg [63:0] mideleg; // @[SIMD_CSR.scala 601:24]
  reg [63:0] mscratch; // @[SIMD_CSR.scala 602:25]
  reg [63:0] pmpcfg0; // @[SIMD_CSR.scala 604:24]
  reg [63:0] pmpcfg1; // @[SIMD_CSR.scala 605:24]
  reg [63:0] pmpcfg2; // @[SIMD_CSR.scala 606:24]
  reg [63:0] pmpcfg3; // @[SIMD_CSR.scala 607:24]
  reg [63:0] pmpaddr0; // @[SIMD_CSR.scala 608:25]
  reg [63:0] pmpaddr1; // @[SIMD_CSR.scala 609:25]
  reg [63:0] pmpaddr2; // @[SIMD_CSR.scala 610:25]
  reg [63:0] pmpaddr3; // @[SIMD_CSR.scala 611:25]
  reg [63:0] vxsat; // @[SIMD_CSR.scala 613:22]
  reg [63:0] stvec; // @[SIMD_CSR.scala 620:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[SIMD_CSR.scala 621:26]
  reg [63:0] satp; // @[SIMD_CSR.scala 623:21]
  reg [63:0] sepc; // @[SIMD_CSR.scala 624:21]
  reg [63:0] scause; // @[SIMD_CSR.scala 625:23]
  reg [63:0] stval; // @[SIMD_CSR.scala 626:18]
  reg [63:0] sscratch; // @[SIMD_CSR.scala 627:25]
  reg [63:0] scounteren; // @[SIMD_CSR.scala 628:27]
  reg [1:0] priviledgeMode; // @[SIMD_CSR.scala 638:31]
  wire [11:0] addr = io_in_bits_src2[16:5]; // @[SIMD_CSR.scala 640:18]
  wire [58:0] _T_29 = io_in_bits_src2[4] ? 59'h7ffffffffffffff : 59'h0; // @[Bitwise.scala 72:12]
  wire [63:0] csri = {_T_29,io_in_bits_src2[4:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_70 = mstatus & 64'h80000003000de122; // @[SIMD_CSR.scala 663:22]
  wire [63:0] _T_103 = mie & sieMask; // @[SIMD_CSR.scala 667:18]
  wire  _T_156 = addr == 12'h302; // @[SIMD_CSR.scala 699:19]
  wire [63:0] _T_205 = vxsat & 64'h1; // @[SIMD_CSR.scala 759:20]
  wire [11:0] _T_208 = {meip,1'h0,meip,1'h0,mtip,1'h0,2'h0,msip,3'h0}; // @[SIMD_CSR.scala 762:22]
  wire [63:0] _GEN_917 = {{52'd0}, _T_208}; // @[SIMD_CSR.scala 762:29]
  wire [63:0] _T_209 = _GEN_917 | mipReg; // @[SIMD_CSR.scala 762:29]
  wire [63:0] _GEN_33 = addr == 12'h344 ? _T_209 : 64'h0; // @[SIMD_CSR.scala 764:29 765:11 768:11]
  wire [63:0] _GEN_36 = addr == 12'h144 ? _T_209 : _GEN_33; // @[SIMD_CSR.scala 761:29 762:11]
  wire [63:0] _GEN_39 = addr == 12'h9 ? _T_205 : _GEN_36; // @[SIMD_CSR.scala 758:31 759:11]
  wire [63:0] _GEN_43 = addr == 12'h3b3 ? pmpaddr3 : _GEN_39; // @[SIMD_CSR.scala 754:43 755:11]
  wire [63:0] _GEN_48 = addr == 12'h3b2 ? pmpaddr2 : _GEN_43; // @[SIMD_CSR.scala 750:43 751:11]
  wire [63:0] _GEN_54 = addr == 12'h3b1 ? pmpaddr1 : _GEN_48; // @[SIMD_CSR.scala 746:43 747:11]
  wire [63:0] _GEN_61 = addr == 12'h3b0 ? pmpaddr0 : _GEN_54; // @[SIMD_CSR.scala 742:43 743:11]
  wire [63:0] _GEN_69 = addr == 12'h3a3 ? pmpcfg3 : _GEN_61; // @[SIMD_CSR.scala 739:33 740:11]
  wire [63:0] _GEN_78 = addr == 12'h3a2 ? pmpcfg2 : _GEN_69; // @[SIMD_CSR.scala 736:33 737:11]
  wire [63:0] _GEN_88 = addr == 12'h3a1 ? pmpcfg1 : _GEN_78; // @[SIMD_CSR.scala 733:33 734:11]
  wire [63:0] _GEN_99 = addr == 12'h3a0 ? pmpcfg0 : _GEN_88; // @[SIMD_CSR.scala 730:33 731:11]
  wire [63:0] _GEN_111 = addr == 12'h343 ? mtval : _GEN_99; // @[SIMD_CSR.scala 727:31 728:11]
  wire [63:0] _GEN_124 = addr == 12'h342 ? mcause : _GEN_111; // @[SIMD_CSR.scala 724:32 725:11]
  wire [63:0] _GEN_138 = addr == 12'h341 ? mepc : _GEN_124; // @[SIMD_CSR.scala 721:30 722:11]
  wire [63:0] _GEN_153 = addr == 12'h340 ? mscratch : _GEN_138; // @[SIMD_CSR.scala 718:34 719:11]
  wire [63:0] _GEN_169 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? 64'h0 : _GEN_153; // @[SIMD_CSR.scala 716:100 717:11]
  wire [63:0] _GEN_185 = addr == 12'h306 ? mcounteren : _GEN_169; // @[SIMD_CSR.scala 713:36 714:11]
  wire [63:0] _GEN_202 = addr == 12'h305 ? mtvec : _GEN_185; // @[SIMD_CSR.scala 710:31 711:11]
  wire [63:0] _GEN_220 = addr == 12'h304 ? mie : _GEN_202; // @[SIMD_CSR.scala 707:29 708:11]
  wire [63:0] _GEN_239 = addr == 12'h303 ? mideleg : _GEN_220; // @[SIMD_CSR.scala 703:33 704:11]
  wire [63:0] _GEN_259 = addr == 12'h302 ? medeleg : _GEN_239; // @[SIMD_CSR.scala 699:33 700:11]
  wire [63:0] _GEN_280 = addr == 12'h301 ? 64'h8000000000141105 : _GEN_259; // @[SIMD_CSR.scala 697:30 698:11]
  wire [63:0] _GEN_301 = addr == 12'h300 ? mstatus : _GEN_280; // @[SIMD_CSR.scala 693:33 694:11]
  wire [63:0] _GEN_323 = addr == 12'h180 ? satp : _GEN_301; // @[SIMD_CSR.scala 687:30 688:11]
  wire [63:0] _GEN_347 = addr == 12'h143 ? stval : _GEN_323; // @[SIMD_CSR.scala 684:31 685:11]
  wire [63:0] _GEN_372 = addr == 12'h142 ? scause : _GEN_347; // @[SIMD_CSR.scala 681:32 682:11]
  wire [63:0] _GEN_398 = addr == 12'h141 ? sepc : _GEN_372; // @[SIMD_CSR.scala 678:30 679:11]
  wire [63:0] _GEN_425 = addr == 12'h140 ? sscratch : _GEN_398; // @[SIMD_CSR.scala 675:34 676:11]
  wire [63:0] _GEN_453 = addr == 12'h106 ? scounteren : _GEN_425; // @[SIMD_CSR.scala 672:36 673:11]
  wire [63:0] _GEN_482 = addr == 12'h105 ? stvec : _GEN_453; // @[SIMD_CSR.scala 669:31 670:11]
  wire [63:0] _GEN_512 = addr == 12'h104 ? _T_103 : _GEN_482; // @[SIMD_CSR.scala 666:29 667:11]
  wire [63:0] rdata = addr == 12'h100 ? _T_70 : _GEN_512; // @[SIMD_CSR.scala 662:27 663:11]
  wire [63:0] _T_30 = rdata | io_in_bits_src1; // @[SIMD_CSR.scala 645:30]
  wire [63:0] _T_31 = ~io_in_bits_src1; // @[SIMD_CSR.scala 646:32]
  wire [63:0] _T_32 = rdata & _T_31; // @[SIMD_CSR.scala 646:30]
  wire [63:0] _T_33 = rdata | csri; // @[SIMD_CSR.scala 648:30]
  wire [63:0] _T_34 = ~csri; // @[SIMD_CSR.scala 649:32]
  wire [63:0] _T_35 = rdata & _T_34; // @[SIMD_CSR.scala 649:30]
  wire  _T_36 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_37 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_38 = 7'h3 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_39 = 7'h5 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_40 = 7'h6 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_41 = 7'h7 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_42 = _T_36 ? io_in_bits_src1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = _T_37 ? _T_30 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = _T_38 ? _T_32 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = _T_39 ? csri : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_40 ? _T_33 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_41 ? _T_35 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_50 = _T_49 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_51 = _T_50 | _T_46; // @[Mux.scala 27:72]
  wire [63:0] wdata = _T_51 | _T_47; // @[Mux.scala 27:72]
  wire  JumpType = io_in_bits_func == 7'h0; // @[SIMD_CSR.scala 653:22]
  wire  _T_55 = ~io_ctrlIn_isMou; // @[SIMD_CSR.scala 654:35]
  wire  wen = io_in_valid & ~JumpType & ~io_ctrlIn_isMou; // @[SIMD_CSR.scala 654:32]
  wire  isIllegalMode = wen & priviledgeMode < addr[9:8]; // @[SIMD_CSR.scala 655:28]
  wire  _T_58 = io_in_bits_func == 7'h2; // @[SIMD_CSR.scala 656:24]
  wire  justRead = (io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6) & io_in_bits_src1 == 64'h0; // @[SIMD_CSR.scala 656:70]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~justRead; // @[SIMD_CSR.scala 657:58]
  wire  RegWen = wen & ~isIllegalWrite & ~isIllegalMode; // @[SIMD_CSR.scala 659:39]
  wire [63:0] _T_72 = mstatus & 64'h39edd; // @[SIMD_CSR.scala 664:24]
  wire [63:0] _T_73 = wdata & 64'hc6122; // @[SIMD_CSR.scala 664:50]
  wire [63:0] _T_74 = _T_72 | _T_73; // @[SIMD_CSR.scala 664:41]
  wire  _T_99 = _T_74[14:13] == 2'h3; // @[SIMD_CSR.scala 665:68]
  wire [63:0] _T_101 = {_T_99,_T_74[62:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_2 = RegWen ? _T_101 : mstatus; // @[SIMD_CSR.scala 665:17 598:24 665:26]
  wire [63:0] _T_106 = ~sieMask; // @[SIMD_CSR.scala 668:64]
  wire [63:0] _T_107 = mie & _T_106; // @[SIMD_CSR.scala 668:62]
  wire [63:0] _T_108 = wdata & sieMask; // @[SIMD_CSR.scala 668:81]
  wire [63:0] _T_109 = _T_107 | _T_108; // @[SIMD_CSR.scala 668:73]
  wire [63:0] _GEN_4 = RegWen ? wdata : stvec; // @[SIMD_CSR.scala 671:17 620:22 671:24]
  wire [63:0] _GEN_5 = RegWen ? wdata : scounteren; // @[SIMD_CSR.scala 674:17 628:27 674:29]
  wire [63:0] _GEN_6 = RegWen ? wdata : sscratch; // @[SIMD_CSR.scala 677:17 627:25 677:27]
  wire [63:0] _GEN_7 = RegWen ? wdata : sepc; // @[SIMD_CSR.scala 680:17 624:21 680:23]
  wire [63:0] _GEN_8 = RegWen ? wdata : scause; // @[SIMD_CSR.scala 683:17 625:23 683:25]
  wire [63:0] _GEN_9 = RegWen ? wdata : stval; // @[SIMD_CSR.scala 686:17 626:18 686:24]
  wire  _T_126 = RegWen & (wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8); // @[SIMD_CSR.scala 689:17]
  wire [63:0] _GEN_10 = RegWen & (wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8) ? wdata : satp; // @[SIMD_CSR.scala 689:113 690:12 623:21]
  wire  _T_152 = wdata[14:13] == 2'h3; // @[SIMD_CSR.scala 696:68]
  wire [63:0] _T_154 = {_T_152,wdata[62:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_12 = RegWen ? _T_154 : mstatus; // @[SIMD_CSR.scala 696:17 598:24 696:26]
  wire [63:0] _T_157 = wdata & 64'hbbff; // @[SIMD_CSR.scala 702:36]
  wire [63:0] _T_159 = medeleg & 64'h4400; // @[SIMD_CSR.scala 702:62]
  wire [63:0] _T_160 = _T_157 | _T_159; // @[SIMD_CSR.scala 702:51]
  wire [63:0] _GEN_13 = RegWen ? _T_160 : medeleg; // @[SIMD_CSR.scala 702:17 600:24 702:26]
  wire [63:0] _T_162 = wdata & 64'h222; // @[SIMD_CSR.scala 706:36]
  wire [63:0] _T_164 = mideleg & 64'h1dd; // @[SIMD_CSR.scala 706:62]
  wire [63:0] _T_165 = _T_162 | _T_164; // @[SIMD_CSR.scala 706:51]
  wire [63:0] _GEN_14 = RegWen ? _T_165 : mideleg; // @[SIMD_CSR.scala 706:17 601:24 706:26]
  wire [63:0] _GEN_15 = RegWen ? wdata : mie; // @[SIMD_CSR.scala 709:17 581:20 709:22]
  wire [63:0] _GEN_16 = RegWen ? wdata : mtvec; // @[SIMD_CSR.scala 712:17 575:22 712:24]
  wire [63:0] _GEN_17 = RegWen ? wdata : mcounteren; // @[SIMD_CSR.scala 715:17 576:27 715:29]
  wire [63:0] _GEN_18 = RegWen ? wdata : mscratch; // @[SIMD_CSR.scala 720:17 602:25 720:27]
  wire [63:0] _GEN_19 = RegWen ? wdata : mepc; // @[SIMD_CSR.scala 579:17 723:{17,23}]
  wire [63:0] _GEN_20 = RegWen ? wdata : mcause; // @[SIMD_CSR.scala 726:17 577:23 726:25]
  wire [63:0] _GEN_21 = RegWen ? wdata : mtval; // @[SIMD_CSR.scala 729:17 578:22 729:24]
  wire [63:0] _GEN_22 = RegWen ? wdata : pmpcfg0; // @[SIMD_CSR.scala 732:17 604:24 732:26]
  wire [63:0] _GEN_23 = RegWen ? wdata : pmpcfg1; // @[SIMD_CSR.scala 735:17 605:24 735:26]
  wire [63:0] _GEN_24 = RegWen ? wdata : pmpcfg2; // @[SIMD_CSR.scala 738:17 606:24 738:26]
  wire [63:0] _GEN_25 = RegWen ? wdata : pmpcfg3; // @[SIMD_CSR.scala 741:17 607:24 741:26]
  wire [63:0] _T_185 = wdata & 64'h3ffffffff; // @[SIMD_CSR.scala 745:37]
  wire [63:0] _GEN_26 = RegWen ? _T_185 : pmpaddr0; // @[SIMD_CSR.scala 745:17 608:25 745:27]
  wire [63:0] _T_190 = wdata & 64'h3fffffc00; // @[SIMD_CSR.scala 749:37]
  wire [63:0] _T_192 = pmpaddr1 & 64'h3ff; // @[SIMD_CSR.scala 749:65]
  wire [63:0] _T_193 = _T_190 | _T_192; // @[SIMD_CSR.scala 749:53]
  wire [63:0] _GEN_27 = RegWen ? _T_193 : pmpaddr1; // @[SIMD_CSR.scala 749:17 609:25 749:27]
  wire [63:0] _T_197 = pmpaddr2 & 64'h3ff; // @[SIMD_CSR.scala 753:65]
  wire [63:0] _T_198 = _T_190 | _T_197; // @[SIMD_CSR.scala 753:53]
  wire [63:0] _GEN_28 = RegWen ? _T_198 : pmpaddr2; // @[SIMD_CSR.scala 753:17 610:25 753:27]
  wire [63:0] _T_202 = pmpaddr3 & 64'h3ff; // @[SIMD_CSR.scala 757:65]
  wire [63:0] _T_203 = _T_190 | _T_202; // @[SIMD_CSR.scala 757:53]
  wire [63:0] _GEN_29 = RegWen ? _T_203 : pmpaddr3; // @[SIMD_CSR.scala 757:17 611:25 757:27]
  wire [63:0] _T_206 = wdata & 64'h1; // @[SIMD_CSR.scala 760:34]
  wire [63:0] _GEN_30 = RegWen ? _T_206 : vxsat; // @[SIMD_CSR.scala 760:17 613:22 760:24]
  wire [63:0] _T_212 = mipReg & _T_106; // @[SIMD_CSR.scala 763:56]
  wire [63:0] _T_213 = _T_108 | _T_212; // @[SIMD_CSR.scala 763:46]
  wire [63:0] _GEN_31 = RegWen ? _T_213 : mipReg; // @[SIMD_CSR.scala 763:17 583:24 763:25]
  wire [63:0] _T_217 = wdata & 64'h77f; // @[SIMD_CSR.scala 766:34]
  wire [63:0] _T_219 = mipReg & 64'h80; // @[SIMD_CSR.scala 766:58]
  wire [63:0] _T_220 = _T_217 | _T_219; // @[SIMD_CSR.scala 766:48]
  wire [63:0] _GEN_32 = RegWen ? _T_220 : mipReg; // @[SIMD_CSR.scala 766:17 583:24 766:24]
  wire [63:0] _GEN_34 = addr == 12'h344 ? _GEN_32 : mipReg; // @[SIMD_CSR.scala 583:24 764:29]
  wire  _GEN_35 = addr == 12'h344 ? 1'h0 : wen; // @[SIMD_CSR.scala 764:29 769:18]
  wire [63:0] _GEN_37 = addr == 12'h144 ? _GEN_31 : _GEN_34; // @[SIMD_CSR.scala 761:29]
  wire  _GEN_38 = addr == 12'h144 ? 1'h0 : _GEN_35; // @[SIMD_CSR.scala 761:29]
  wire [63:0] _GEN_40 = addr == 12'h9 ? _GEN_30 : vxsat; // @[SIMD_CSR.scala 613:22 758:31]
  wire [63:0] _GEN_41 = addr == 12'h9 ? mipReg : _GEN_37; // @[SIMD_CSR.scala 583:24 758:31]
  wire  _GEN_42 = addr == 12'h9 ? 1'h0 : _GEN_38; // @[SIMD_CSR.scala 758:31]
  wire [63:0] _GEN_44 = addr == 12'h3b3 ? _GEN_29 : pmpaddr3; // @[SIMD_CSR.scala 611:25 754:43]
  wire [63:0] _GEN_45 = addr == 12'h3b3 ? vxsat : _GEN_40; // @[SIMD_CSR.scala 613:22 754:43]
  wire [63:0] _GEN_46 = addr == 12'h3b3 ? mipReg : _GEN_41; // @[SIMD_CSR.scala 583:24 754:43]
  wire  _GEN_47 = addr == 12'h3b3 ? 1'h0 : _GEN_42; // @[SIMD_CSR.scala 754:43]
  wire [63:0] _GEN_49 = addr == 12'h3b2 ? _GEN_28 : pmpaddr2; // @[SIMD_CSR.scala 610:25 750:43]
  wire [63:0] _GEN_50 = addr == 12'h3b2 ? pmpaddr3 : _GEN_44; // @[SIMD_CSR.scala 611:25 750:43]
  wire [63:0] _GEN_51 = addr == 12'h3b2 ? vxsat : _GEN_45; // @[SIMD_CSR.scala 613:22 750:43]
  wire [63:0] _GEN_52 = addr == 12'h3b2 ? mipReg : _GEN_46; // @[SIMD_CSR.scala 583:24 750:43]
  wire  _GEN_53 = addr == 12'h3b2 ? 1'h0 : _GEN_47; // @[SIMD_CSR.scala 750:43]
  wire [63:0] _GEN_55 = addr == 12'h3b1 ? _GEN_27 : pmpaddr1; // @[SIMD_CSR.scala 609:25 746:43]
  wire [63:0] _GEN_56 = addr == 12'h3b1 ? pmpaddr2 : _GEN_49; // @[SIMD_CSR.scala 610:25 746:43]
  wire [63:0] _GEN_57 = addr == 12'h3b1 ? pmpaddr3 : _GEN_50; // @[SIMD_CSR.scala 611:25 746:43]
  wire [63:0] _GEN_58 = addr == 12'h3b1 ? vxsat : _GEN_51; // @[SIMD_CSR.scala 613:22 746:43]
  wire [63:0] _GEN_59 = addr == 12'h3b1 ? mipReg : _GEN_52; // @[SIMD_CSR.scala 583:24 746:43]
  wire  _GEN_60 = addr == 12'h3b1 ? 1'h0 : _GEN_53; // @[SIMD_CSR.scala 746:43]
  wire [63:0] _GEN_62 = addr == 12'h3b0 ? _GEN_26 : pmpaddr0; // @[SIMD_CSR.scala 608:25 742:43]
  wire [63:0] _GEN_63 = addr == 12'h3b0 ? pmpaddr1 : _GEN_55; // @[SIMD_CSR.scala 609:25 742:43]
  wire [63:0] _GEN_64 = addr == 12'h3b0 ? pmpaddr2 : _GEN_56; // @[SIMD_CSR.scala 610:25 742:43]
  wire [63:0] _GEN_65 = addr == 12'h3b0 ? pmpaddr3 : _GEN_57; // @[SIMD_CSR.scala 611:25 742:43]
  wire [63:0] _GEN_66 = addr == 12'h3b0 ? vxsat : _GEN_58; // @[SIMD_CSR.scala 613:22 742:43]
  wire [63:0] _GEN_67 = addr == 12'h3b0 ? mipReg : _GEN_59; // @[SIMD_CSR.scala 583:24 742:43]
  wire  _GEN_68 = addr == 12'h3b0 ? 1'h0 : _GEN_60; // @[SIMD_CSR.scala 742:43]
  wire [63:0] _GEN_70 = addr == 12'h3a3 ? _GEN_25 : pmpcfg3; // @[SIMD_CSR.scala 607:24 739:33]
  wire [63:0] _GEN_71 = addr == 12'h3a3 ? pmpaddr0 : _GEN_62; // @[SIMD_CSR.scala 608:25 739:33]
  wire [63:0] _GEN_72 = addr == 12'h3a3 ? pmpaddr1 : _GEN_63; // @[SIMD_CSR.scala 609:25 739:33]
  wire [63:0] _GEN_73 = addr == 12'h3a3 ? pmpaddr2 : _GEN_64; // @[SIMD_CSR.scala 610:25 739:33]
  wire [63:0] _GEN_74 = addr == 12'h3a3 ? pmpaddr3 : _GEN_65; // @[SIMD_CSR.scala 611:25 739:33]
  wire [63:0] _GEN_75 = addr == 12'h3a3 ? vxsat : _GEN_66; // @[SIMD_CSR.scala 613:22 739:33]
  wire [63:0] _GEN_76 = addr == 12'h3a3 ? mipReg : _GEN_67; // @[SIMD_CSR.scala 583:24 739:33]
  wire  _GEN_77 = addr == 12'h3a3 ? 1'h0 : _GEN_68; // @[SIMD_CSR.scala 739:33]
  wire [63:0] _GEN_79 = addr == 12'h3a2 ? _GEN_24 : pmpcfg2; // @[SIMD_CSR.scala 606:24 736:33]
  wire [63:0] _GEN_80 = addr == 12'h3a2 ? pmpcfg3 : _GEN_70; // @[SIMD_CSR.scala 607:24 736:33]
  wire [63:0] _GEN_81 = addr == 12'h3a2 ? pmpaddr0 : _GEN_71; // @[SIMD_CSR.scala 608:25 736:33]
  wire [63:0] _GEN_82 = addr == 12'h3a2 ? pmpaddr1 : _GEN_72; // @[SIMD_CSR.scala 609:25 736:33]
  wire [63:0] _GEN_83 = addr == 12'h3a2 ? pmpaddr2 : _GEN_73; // @[SIMD_CSR.scala 610:25 736:33]
  wire [63:0] _GEN_84 = addr == 12'h3a2 ? pmpaddr3 : _GEN_74; // @[SIMD_CSR.scala 611:25 736:33]
  wire [63:0] _GEN_85 = addr == 12'h3a2 ? vxsat : _GEN_75; // @[SIMD_CSR.scala 613:22 736:33]
  wire [63:0] _GEN_86 = addr == 12'h3a2 ? mipReg : _GEN_76; // @[SIMD_CSR.scala 583:24 736:33]
  wire  _GEN_87 = addr == 12'h3a2 ? 1'h0 : _GEN_77; // @[SIMD_CSR.scala 736:33]
  wire [63:0] _GEN_89 = addr == 12'h3a1 ? _GEN_23 : pmpcfg1; // @[SIMD_CSR.scala 605:24 733:33]
  wire [63:0] _GEN_90 = addr == 12'h3a1 ? pmpcfg2 : _GEN_79; // @[SIMD_CSR.scala 606:24 733:33]
  wire [63:0] _GEN_91 = addr == 12'h3a1 ? pmpcfg3 : _GEN_80; // @[SIMD_CSR.scala 607:24 733:33]
  wire [63:0] _GEN_92 = addr == 12'h3a1 ? pmpaddr0 : _GEN_81; // @[SIMD_CSR.scala 608:25 733:33]
  wire [63:0] _GEN_93 = addr == 12'h3a1 ? pmpaddr1 : _GEN_82; // @[SIMD_CSR.scala 609:25 733:33]
  wire [63:0] _GEN_94 = addr == 12'h3a1 ? pmpaddr2 : _GEN_83; // @[SIMD_CSR.scala 610:25 733:33]
  wire [63:0] _GEN_95 = addr == 12'h3a1 ? pmpaddr3 : _GEN_84; // @[SIMD_CSR.scala 611:25 733:33]
  wire [63:0] _GEN_96 = addr == 12'h3a1 ? vxsat : _GEN_85; // @[SIMD_CSR.scala 613:22 733:33]
  wire [63:0] _GEN_97 = addr == 12'h3a1 ? mipReg : _GEN_86; // @[SIMD_CSR.scala 583:24 733:33]
  wire  _GEN_98 = addr == 12'h3a1 ? 1'h0 : _GEN_87; // @[SIMD_CSR.scala 733:33]
  wire [63:0] _GEN_100 = addr == 12'h3a0 ? _GEN_22 : pmpcfg0; // @[SIMD_CSR.scala 604:24 730:33]
  wire [63:0] _GEN_101 = addr == 12'h3a0 ? pmpcfg1 : _GEN_89; // @[SIMD_CSR.scala 605:24 730:33]
  wire [63:0] _GEN_102 = addr == 12'h3a0 ? pmpcfg2 : _GEN_90; // @[SIMD_CSR.scala 606:24 730:33]
  wire [63:0] _GEN_103 = addr == 12'h3a0 ? pmpcfg3 : _GEN_91; // @[SIMD_CSR.scala 607:24 730:33]
  wire [63:0] _GEN_104 = addr == 12'h3a0 ? pmpaddr0 : _GEN_92; // @[SIMD_CSR.scala 608:25 730:33]
  wire [63:0] _GEN_105 = addr == 12'h3a0 ? pmpaddr1 : _GEN_93; // @[SIMD_CSR.scala 609:25 730:33]
  wire [63:0] _GEN_106 = addr == 12'h3a0 ? pmpaddr2 : _GEN_94; // @[SIMD_CSR.scala 610:25 730:33]
  wire [63:0] _GEN_107 = addr == 12'h3a0 ? pmpaddr3 : _GEN_95; // @[SIMD_CSR.scala 611:25 730:33]
  wire [63:0] _GEN_108 = addr == 12'h3a0 ? vxsat : _GEN_96; // @[SIMD_CSR.scala 613:22 730:33]
  wire [63:0] _GEN_109 = addr == 12'h3a0 ? mipReg : _GEN_97; // @[SIMD_CSR.scala 583:24 730:33]
  wire  _GEN_110 = addr == 12'h3a0 ? 1'h0 : _GEN_98; // @[SIMD_CSR.scala 730:33]
  wire [63:0] _GEN_112 = addr == 12'h343 ? _GEN_21 : mtval; // @[SIMD_CSR.scala 578:22 727:31]
  wire [63:0] _GEN_113 = addr == 12'h343 ? pmpcfg0 : _GEN_100; // @[SIMD_CSR.scala 604:24 727:31]
  wire [63:0] _GEN_114 = addr == 12'h343 ? pmpcfg1 : _GEN_101; // @[SIMD_CSR.scala 605:24 727:31]
  wire [63:0] _GEN_115 = addr == 12'h343 ? pmpcfg2 : _GEN_102; // @[SIMD_CSR.scala 606:24 727:31]
  wire [63:0] _GEN_116 = addr == 12'h343 ? pmpcfg3 : _GEN_103; // @[SIMD_CSR.scala 607:24 727:31]
  wire [63:0] _GEN_117 = addr == 12'h343 ? pmpaddr0 : _GEN_104; // @[SIMD_CSR.scala 608:25 727:31]
  wire [63:0] _GEN_118 = addr == 12'h343 ? pmpaddr1 : _GEN_105; // @[SIMD_CSR.scala 609:25 727:31]
  wire [63:0] _GEN_119 = addr == 12'h343 ? pmpaddr2 : _GEN_106; // @[SIMD_CSR.scala 610:25 727:31]
  wire [63:0] _GEN_120 = addr == 12'h343 ? pmpaddr3 : _GEN_107; // @[SIMD_CSR.scala 611:25 727:31]
  wire [63:0] _GEN_121 = addr == 12'h343 ? vxsat : _GEN_108; // @[SIMD_CSR.scala 613:22 727:31]
  wire [63:0] _GEN_122 = addr == 12'h343 ? mipReg : _GEN_109; // @[SIMD_CSR.scala 583:24 727:31]
  wire  _GEN_123 = addr == 12'h343 ? 1'h0 : _GEN_110; // @[SIMD_CSR.scala 727:31]
  wire [63:0] _GEN_125 = addr == 12'h342 ? _GEN_20 : mcause; // @[SIMD_CSR.scala 577:23 724:32]
  wire [63:0] _GEN_126 = addr == 12'h342 ? mtval : _GEN_112; // @[SIMD_CSR.scala 578:22 724:32]
  wire [63:0] _GEN_127 = addr == 12'h342 ? pmpcfg0 : _GEN_113; // @[SIMD_CSR.scala 604:24 724:32]
  wire [63:0] _GEN_128 = addr == 12'h342 ? pmpcfg1 : _GEN_114; // @[SIMD_CSR.scala 605:24 724:32]
  wire [63:0] _GEN_129 = addr == 12'h342 ? pmpcfg2 : _GEN_115; // @[SIMD_CSR.scala 606:24 724:32]
  wire [63:0] _GEN_130 = addr == 12'h342 ? pmpcfg3 : _GEN_116; // @[SIMD_CSR.scala 607:24 724:32]
  wire [63:0] _GEN_131 = addr == 12'h342 ? pmpaddr0 : _GEN_117; // @[SIMD_CSR.scala 608:25 724:32]
  wire [63:0] _GEN_132 = addr == 12'h342 ? pmpaddr1 : _GEN_118; // @[SIMD_CSR.scala 609:25 724:32]
  wire [63:0] _GEN_133 = addr == 12'h342 ? pmpaddr2 : _GEN_119; // @[SIMD_CSR.scala 610:25 724:32]
  wire [63:0] _GEN_134 = addr == 12'h342 ? pmpaddr3 : _GEN_120; // @[SIMD_CSR.scala 611:25 724:32]
  wire [63:0] _GEN_135 = addr == 12'h342 ? vxsat : _GEN_121; // @[SIMD_CSR.scala 613:22 724:32]
  wire [63:0] _GEN_136 = addr == 12'h342 ? mipReg : _GEN_122; // @[SIMD_CSR.scala 583:24 724:32]
  wire  _GEN_137 = addr == 12'h342 ? 1'h0 : _GEN_123; // @[SIMD_CSR.scala 724:32]
  wire [63:0] _GEN_139 = addr == 12'h341 ? _GEN_19 : mepc; // @[SIMD_CSR.scala 579:17 721:30]
  wire [63:0] _GEN_140 = addr == 12'h341 ? mcause : _GEN_125; // @[SIMD_CSR.scala 577:23 721:30]
  wire [63:0] _GEN_141 = addr == 12'h341 ? mtval : _GEN_126; // @[SIMD_CSR.scala 578:22 721:30]
  wire [63:0] _GEN_142 = addr == 12'h341 ? pmpcfg0 : _GEN_127; // @[SIMD_CSR.scala 604:24 721:30]
  wire [63:0] _GEN_143 = addr == 12'h341 ? pmpcfg1 : _GEN_128; // @[SIMD_CSR.scala 605:24 721:30]
  wire [63:0] _GEN_144 = addr == 12'h341 ? pmpcfg2 : _GEN_129; // @[SIMD_CSR.scala 606:24 721:30]
  wire [63:0] _GEN_145 = addr == 12'h341 ? pmpcfg3 : _GEN_130; // @[SIMD_CSR.scala 607:24 721:30]
  wire [63:0] _GEN_146 = addr == 12'h341 ? pmpaddr0 : _GEN_131; // @[SIMD_CSR.scala 608:25 721:30]
  wire [63:0] _GEN_147 = addr == 12'h341 ? pmpaddr1 : _GEN_132; // @[SIMD_CSR.scala 609:25 721:30]
  wire [63:0] _GEN_148 = addr == 12'h341 ? pmpaddr2 : _GEN_133; // @[SIMD_CSR.scala 610:25 721:30]
  wire [63:0] _GEN_149 = addr == 12'h341 ? pmpaddr3 : _GEN_134; // @[SIMD_CSR.scala 611:25 721:30]
  wire [63:0] _GEN_150 = addr == 12'h341 ? vxsat : _GEN_135; // @[SIMD_CSR.scala 613:22 721:30]
  wire [63:0] _GEN_151 = addr == 12'h341 ? mipReg : _GEN_136; // @[SIMD_CSR.scala 583:24 721:30]
  wire  _GEN_152 = addr == 12'h341 ? 1'h0 : _GEN_137; // @[SIMD_CSR.scala 721:30]
  wire [63:0] _GEN_154 = addr == 12'h340 ? _GEN_18 : mscratch; // @[SIMD_CSR.scala 602:25 718:34]
  wire [63:0] _GEN_155 = addr == 12'h340 ? mepc : _GEN_139; // @[SIMD_CSR.scala 579:17 718:34]
  wire [63:0] _GEN_156 = addr == 12'h340 ? mcause : _GEN_140; // @[SIMD_CSR.scala 577:23 718:34]
  wire [63:0] _GEN_157 = addr == 12'h340 ? mtval : _GEN_141; // @[SIMD_CSR.scala 578:22 718:34]
  wire [63:0] _GEN_158 = addr == 12'h340 ? pmpcfg0 : _GEN_142; // @[SIMD_CSR.scala 604:24 718:34]
  wire [63:0] _GEN_159 = addr == 12'h340 ? pmpcfg1 : _GEN_143; // @[SIMD_CSR.scala 605:24 718:34]
  wire [63:0] _GEN_160 = addr == 12'h340 ? pmpcfg2 : _GEN_144; // @[SIMD_CSR.scala 606:24 718:34]
  wire [63:0] _GEN_161 = addr == 12'h340 ? pmpcfg3 : _GEN_145; // @[SIMD_CSR.scala 607:24 718:34]
  wire [63:0] _GEN_162 = addr == 12'h340 ? pmpaddr0 : _GEN_146; // @[SIMD_CSR.scala 608:25 718:34]
  wire [63:0] _GEN_163 = addr == 12'h340 ? pmpaddr1 : _GEN_147; // @[SIMD_CSR.scala 609:25 718:34]
  wire [63:0] _GEN_164 = addr == 12'h340 ? pmpaddr2 : _GEN_148; // @[SIMD_CSR.scala 610:25 718:34]
  wire [63:0] _GEN_165 = addr == 12'h340 ? pmpaddr3 : _GEN_149; // @[SIMD_CSR.scala 611:25 718:34]
  wire [63:0] _GEN_166 = addr == 12'h340 ? vxsat : _GEN_150; // @[SIMD_CSR.scala 613:22 718:34]
  wire [63:0] _GEN_167 = addr == 12'h340 ? mipReg : _GEN_151; // @[SIMD_CSR.scala 583:24 718:34]
  wire  _GEN_168 = addr == 12'h340 ? 1'h0 : _GEN_152; // @[SIMD_CSR.scala 718:34]
  wire [63:0] _GEN_170 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? mscratch : _GEN_154; // @[SIMD_CSR.scala 716:100 602:25]
  wire [63:0] _GEN_171 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? mepc : _GEN_155; // @[SIMD_CSR.scala 716:100 579:17]
  wire [63:0] _GEN_172 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? mcause : _GEN_156; // @[SIMD_CSR.scala 716:100 577:23]
  wire [63:0] _GEN_173 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? mtval : _GEN_157; // @[SIMD_CSR.scala 716:100 578:22]
  wire [63:0] _GEN_174 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpcfg0 : _GEN_158; // @[SIMD_CSR.scala 716:100 604:24]
  wire [63:0] _GEN_175 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpcfg1 : _GEN_159; // @[SIMD_CSR.scala 716:100 605:24]
  wire [63:0] _GEN_176 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpcfg2 : _GEN_160; // @[SIMD_CSR.scala 716:100 606:24]
  wire [63:0] _GEN_177 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpcfg3 : _GEN_161; // @[SIMD_CSR.scala 716:100 607:24]
  wire [63:0] _GEN_178 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpaddr0 : _GEN_162; // @[SIMD_CSR.scala 716:100 608:25]
  wire [63:0] _GEN_179 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpaddr1 : _GEN_163; // @[SIMD_CSR.scala 716:100 609:25]
  wire [63:0] _GEN_180 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpaddr2 : _GEN_164; // @[SIMD_CSR.scala 716:100 610:25]
  wire [63:0] _GEN_181 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? pmpaddr3 : _GEN_165; // @[SIMD_CSR.scala 716:100 611:25]
  wire [63:0] _GEN_182 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? vxsat : _GEN_166; // @[SIMD_CSR.scala 716:100 613:22]
  wire [63:0] _GEN_183 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? mipReg : _GEN_167; // @[SIMD_CSR.scala 716:100 583:24]
  wire  _GEN_184 = addr == 12'hf11 | addr == 12'hf12 | addr == 12'hf13 | addr == 12'hf14 ? 1'h0 : _GEN_168; // @[SIMD_CSR.scala 716:100]
  wire [63:0] _GEN_186 = addr == 12'h306 ? _GEN_17 : mcounteren; // @[SIMD_CSR.scala 576:27 713:36]
  wire [63:0] _GEN_187 = addr == 12'h306 ? mscratch : _GEN_170; // @[SIMD_CSR.scala 602:25 713:36]
  wire [63:0] _GEN_188 = addr == 12'h306 ? mepc : _GEN_171; // @[SIMD_CSR.scala 579:17 713:36]
  wire [63:0] _GEN_189 = addr == 12'h306 ? mcause : _GEN_172; // @[SIMD_CSR.scala 577:23 713:36]
  wire [63:0] _GEN_190 = addr == 12'h306 ? mtval : _GEN_173; // @[SIMD_CSR.scala 578:22 713:36]
  wire [63:0] _GEN_191 = addr == 12'h306 ? pmpcfg0 : _GEN_174; // @[SIMD_CSR.scala 604:24 713:36]
  wire [63:0] _GEN_192 = addr == 12'h306 ? pmpcfg1 : _GEN_175; // @[SIMD_CSR.scala 605:24 713:36]
  wire [63:0] _GEN_193 = addr == 12'h306 ? pmpcfg2 : _GEN_176; // @[SIMD_CSR.scala 606:24 713:36]
  wire [63:0] _GEN_194 = addr == 12'h306 ? pmpcfg3 : _GEN_177; // @[SIMD_CSR.scala 607:24 713:36]
  wire [63:0] _GEN_195 = addr == 12'h306 ? pmpaddr0 : _GEN_178; // @[SIMD_CSR.scala 608:25 713:36]
  wire [63:0] _GEN_196 = addr == 12'h306 ? pmpaddr1 : _GEN_179; // @[SIMD_CSR.scala 609:25 713:36]
  wire [63:0] _GEN_197 = addr == 12'h306 ? pmpaddr2 : _GEN_180; // @[SIMD_CSR.scala 610:25 713:36]
  wire [63:0] _GEN_198 = addr == 12'h306 ? pmpaddr3 : _GEN_181; // @[SIMD_CSR.scala 611:25 713:36]
  wire [63:0] _GEN_199 = addr == 12'h306 ? vxsat : _GEN_182; // @[SIMD_CSR.scala 613:22 713:36]
  wire [63:0] _GEN_200 = addr == 12'h306 ? mipReg : _GEN_183; // @[SIMD_CSR.scala 583:24 713:36]
  wire  _GEN_201 = addr == 12'h306 ? 1'h0 : _GEN_184; // @[SIMD_CSR.scala 713:36]
  wire [63:0] _GEN_203 = addr == 12'h305 ? _GEN_16 : mtvec; // @[SIMD_CSR.scala 575:22 710:31]
  wire [63:0] _GEN_204 = addr == 12'h305 ? mcounteren : _GEN_186; // @[SIMD_CSR.scala 576:27 710:31]
  wire [63:0] _GEN_205 = addr == 12'h305 ? mscratch : _GEN_187; // @[SIMD_CSR.scala 602:25 710:31]
  wire [63:0] _GEN_206 = addr == 12'h305 ? mepc : _GEN_188; // @[SIMD_CSR.scala 579:17 710:31]
  wire [63:0] _GEN_207 = addr == 12'h305 ? mcause : _GEN_189; // @[SIMD_CSR.scala 577:23 710:31]
  wire [63:0] _GEN_208 = addr == 12'h305 ? mtval : _GEN_190; // @[SIMD_CSR.scala 578:22 710:31]
  wire [63:0] _GEN_209 = addr == 12'h305 ? pmpcfg0 : _GEN_191; // @[SIMD_CSR.scala 604:24 710:31]
  wire [63:0] _GEN_210 = addr == 12'h305 ? pmpcfg1 : _GEN_192; // @[SIMD_CSR.scala 605:24 710:31]
  wire [63:0] _GEN_211 = addr == 12'h305 ? pmpcfg2 : _GEN_193; // @[SIMD_CSR.scala 606:24 710:31]
  wire [63:0] _GEN_212 = addr == 12'h305 ? pmpcfg3 : _GEN_194; // @[SIMD_CSR.scala 607:24 710:31]
  wire [63:0] _GEN_213 = addr == 12'h305 ? pmpaddr0 : _GEN_195; // @[SIMD_CSR.scala 608:25 710:31]
  wire [63:0] _GEN_214 = addr == 12'h305 ? pmpaddr1 : _GEN_196; // @[SIMD_CSR.scala 609:25 710:31]
  wire [63:0] _GEN_215 = addr == 12'h305 ? pmpaddr2 : _GEN_197; // @[SIMD_CSR.scala 610:25 710:31]
  wire [63:0] _GEN_216 = addr == 12'h305 ? pmpaddr3 : _GEN_198; // @[SIMD_CSR.scala 611:25 710:31]
  wire [63:0] _GEN_217 = addr == 12'h305 ? vxsat : _GEN_199; // @[SIMD_CSR.scala 613:22 710:31]
  wire [63:0] _GEN_218 = addr == 12'h305 ? mipReg : _GEN_200; // @[SIMD_CSR.scala 583:24 710:31]
  wire  _GEN_219 = addr == 12'h305 ? 1'h0 : _GEN_201; // @[SIMD_CSR.scala 710:31]
  wire [63:0] _GEN_221 = addr == 12'h304 ? _GEN_15 : mie; // @[SIMD_CSR.scala 581:20 707:29]
  wire [63:0] _GEN_222 = addr == 12'h304 ? mtvec : _GEN_203; // @[SIMD_CSR.scala 575:22 707:29]
  wire [63:0] _GEN_223 = addr == 12'h304 ? mcounteren : _GEN_204; // @[SIMD_CSR.scala 576:27 707:29]
  wire [63:0] _GEN_224 = addr == 12'h304 ? mscratch : _GEN_205; // @[SIMD_CSR.scala 602:25 707:29]
  wire [63:0] _GEN_225 = addr == 12'h304 ? mepc : _GEN_206; // @[SIMD_CSR.scala 579:17 707:29]
  wire [63:0] _GEN_226 = addr == 12'h304 ? mcause : _GEN_207; // @[SIMD_CSR.scala 577:23 707:29]
  wire [63:0] _GEN_227 = addr == 12'h304 ? mtval : _GEN_208; // @[SIMD_CSR.scala 578:22 707:29]
  wire [63:0] _GEN_228 = addr == 12'h304 ? pmpcfg0 : _GEN_209; // @[SIMD_CSR.scala 604:24 707:29]
  wire [63:0] _GEN_229 = addr == 12'h304 ? pmpcfg1 : _GEN_210; // @[SIMD_CSR.scala 605:24 707:29]
  wire [63:0] _GEN_230 = addr == 12'h304 ? pmpcfg2 : _GEN_211; // @[SIMD_CSR.scala 606:24 707:29]
  wire [63:0] _GEN_231 = addr == 12'h304 ? pmpcfg3 : _GEN_212; // @[SIMD_CSR.scala 607:24 707:29]
  wire [63:0] _GEN_232 = addr == 12'h304 ? pmpaddr0 : _GEN_213; // @[SIMD_CSR.scala 608:25 707:29]
  wire [63:0] _GEN_233 = addr == 12'h304 ? pmpaddr1 : _GEN_214; // @[SIMD_CSR.scala 609:25 707:29]
  wire [63:0] _GEN_234 = addr == 12'h304 ? pmpaddr2 : _GEN_215; // @[SIMD_CSR.scala 610:25 707:29]
  wire [63:0] _GEN_235 = addr == 12'h304 ? pmpaddr3 : _GEN_216; // @[SIMD_CSR.scala 611:25 707:29]
  wire [63:0] _GEN_236 = addr == 12'h304 ? vxsat : _GEN_217; // @[SIMD_CSR.scala 613:22 707:29]
  wire [63:0] _GEN_237 = addr == 12'h304 ? mipReg : _GEN_218; // @[SIMD_CSR.scala 583:24 707:29]
  wire  _GEN_238 = addr == 12'h304 ? 1'h0 : _GEN_219; // @[SIMD_CSR.scala 707:29]
  wire [63:0] _GEN_240 = addr == 12'h303 ? _GEN_14 : mideleg; // @[SIMD_CSR.scala 601:24 703:33]
  wire [63:0] _GEN_241 = addr == 12'h303 ? mie : _GEN_221; // @[SIMD_CSR.scala 581:20 703:33]
  wire [63:0] _GEN_242 = addr == 12'h303 ? mtvec : _GEN_222; // @[SIMD_CSR.scala 575:22 703:33]
  wire [63:0] _GEN_243 = addr == 12'h303 ? mcounteren : _GEN_223; // @[SIMD_CSR.scala 576:27 703:33]
  wire [63:0] _GEN_244 = addr == 12'h303 ? mscratch : _GEN_224; // @[SIMD_CSR.scala 602:25 703:33]
  wire [63:0] _GEN_245 = addr == 12'h303 ? mepc : _GEN_225; // @[SIMD_CSR.scala 579:17 703:33]
  wire [63:0] _GEN_246 = addr == 12'h303 ? mcause : _GEN_226; // @[SIMD_CSR.scala 577:23 703:33]
  wire [63:0] _GEN_247 = addr == 12'h303 ? mtval : _GEN_227; // @[SIMD_CSR.scala 578:22 703:33]
  wire [63:0] _GEN_248 = addr == 12'h303 ? pmpcfg0 : _GEN_228; // @[SIMD_CSR.scala 604:24 703:33]
  wire [63:0] _GEN_249 = addr == 12'h303 ? pmpcfg1 : _GEN_229; // @[SIMD_CSR.scala 605:24 703:33]
  wire [63:0] _GEN_250 = addr == 12'h303 ? pmpcfg2 : _GEN_230; // @[SIMD_CSR.scala 606:24 703:33]
  wire [63:0] _GEN_251 = addr == 12'h303 ? pmpcfg3 : _GEN_231; // @[SIMD_CSR.scala 607:24 703:33]
  wire [63:0] _GEN_252 = addr == 12'h303 ? pmpaddr0 : _GEN_232; // @[SIMD_CSR.scala 608:25 703:33]
  wire [63:0] _GEN_253 = addr == 12'h303 ? pmpaddr1 : _GEN_233; // @[SIMD_CSR.scala 609:25 703:33]
  wire [63:0] _GEN_254 = addr == 12'h303 ? pmpaddr2 : _GEN_234; // @[SIMD_CSR.scala 610:25 703:33]
  wire [63:0] _GEN_255 = addr == 12'h303 ? pmpaddr3 : _GEN_235; // @[SIMD_CSR.scala 611:25 703:33]
  wire [63:0] _GEN_256 = addr == 12'h303 ? vxsat : _GEN_236; // @[SIMD_CSR.scala 613:22 703:33]
  wire [63:0] _GEN_257 = addr == 12'h303 ? mipReg : _GEN_237; // @[SIMD_CSR.scala 583:24 703:33]
  wire  _GEN_258 = addr == 12'h303 ? 1'h0 : _GEN_238; // @[SIMD_CSR.scala 703:33]
  wire [63:0] _GEN_260 = addr == 12'h302 ? _GEN_13 : medeleg; // @[SIMD_CSR.scala 600:24 699:33]
  wire [63:0] _GEN_261 = addr == 12'h302 ? mideleg : _GEN_240; // @[SIMD_CSR.scala 601:24 699:33]
  wire [63:0] _GEN_262 = addr == 12'h302 ? mie : _GEN_241; // @[SIMD_CSR.scala 581:20 699:33]
  wire [63:0] _GEN_263 = addr == 12'h302 ? mtvec : _GEN_242; // @[SIMD_CSR.scala 575:22 699:33]
  wire [63:0] _GEN_264 = addr == 12'h302 ? mcounteren : _GEN_243; // @[SIMD_CSR.scala 576:27 699:33]
  wire [63:0] _GEN_265 = addr == 12'h302 ? mscratch : _GEN_244; // @[SIMD_CSR.scala 602:25 699:33]
  wire [63:0] _GEN_266 = addr == 12'h302 ? mepc : _GEN_245; // @[SIMD_CSR.scala 579:17 699:33]
  wire [63:0] _GEN_267 = addr == 12'h302 ? mcause : _GEN_246; // @[SIMD_CSR.scala 577:23 699:33]
  wire [63:0] _GEN_268 = addr == 12'h302 ? mtval : _GEN_247; // @[SIMD_CSR.scala 578:22 699:33]
  wire [63:0] _GEN_269 = addr == 12'h302 ? pmpcfg0 : _GEN_248; // @[SIMD_CSR.scala 604:24 699:33]
  wire [63:0] _GEN_270 = addr == 12'h302 ? pmpcfg1 : _GEN_249; // @[SIMD_CSR.scala 605:24 699:33]
  wire [63:0] _GEN_271 = addr == 12'h302 ? pmpcfg2 : _GEN_250; // @[SIMD_CSR.scala 606:24 699:33]
  wire [63:0] _GEN_272 = addr == 12'h302 ? pmpcfg3 : _GEN_251; // @[SIMD_CSR.scala 607:24 699:33]
  wire [63:0] _GEN_273 = addr == 12'h302 ? pmpaddr0 : _GEN_252; // @[SIMD_CSR.scala 608:25 699:33]
  wire [63:0] _GEN_274 = addr == 12'h302 ? pmpaddr1 : _GEN_253; // @[SIMD_CSR.scala 609:25 699:33]
  wire [63:0] _GEN_275 = addr == 12'h302 ? pmpaddr2 : _GEN_254; // @[SIMD_CSR.scala 610:25 699:33]
  wire [63:0] _GEN_276 = addr == 12'h302 ? pmpaddr3 : _GEN_255; // @[SIMD_CSR.scala 611:25 699:33]
  wire [63:0] _GEN_277 = addr == 12'h302 ? vxsat : _GEN_256; // @[SIMD_CSR.scala 613:22 699:33]
  wire [63:0] _GEN_278 = addr == 12'h302 ? mipReg : _GEN_257; // @[SIMD_CSR.scala 583:24 699:33]
  wire  _GEN_279 = addr == 12'h302 ? 1'h0 : _GEN_258; // @[SIMD_CSR.scala 699:33]
  wire [63:0] _GEN_281 = addr == 12'h301 ? medeleg : _GEN_260; // @[SIMD_CSR.scala 600:24 697:30]
  wire [63:0] _GEN_282 = addr == 12'h301 ? mideleg : _GEN_261; // @[SIMD_CSR.scala 601:24 697:30]
  wire [63:0] _GEN_283 = addr == 12'h301 ? mie : _GEN_262; // @[SIMD_CSR.scala 581:20 697:30]
  wire [63:0] _GEN_284 = addr == 12'h301 ? mtvec : _GEN_263; // @[SIMD_CSR.scala 575:22 697:30]
  wire [63:0] _GEN_285 = addr == 12'h301 ? mcounteren : _GEN_264; // @[SIMD_CSR.scala 576:27 697:30]
  wire [63:0] _GEN_286 = addr == 12'h301 ? mscratch : _GEN_265; // @[SIMD_CSR.scala 602:25 697:30]
  wire [63:0] _GEN_287 = addr == 12'h301 ? mepc : _GEN_266; // @[SIMD_CSR.scala 579:17 697:30]
  wire [63:0] _GEN_288 = addr == 12'h301 ? mcause : _GEN_267; // @[SIMD_CSR.scala 577:23 697:30]
  wire [63:0] _GEN_289 = addr == 12'h301 ? mtval : _GEN_268; // @[SIMD_CSR.scala 578:22 697:30]
  wire [63:0] _GEN_290 = addr == 12'h301 ? pmpcfg0 : _GEN_269; // @[SIMD_CSR.scala 604:24 697:30]
  wire [63:0] _GEN_291 = addr == 12'h301 ? pmpcfg1 : _GEN_270; // @[SIMD_CSR.scala 605:24 697:30]
  wire [63:0] _GEN_292 = addr == 12'h301 ? pmpcfg2 : _GEN_271; // @[SIMD_CSR.scala 606:24 697:30]
  wire [63:0] _GEN_293 = addr == 12'h301 ? pmpcfg3 : _GEN_272; // @[SIMD_CSR.scala 607:24 697:30]
  wire [63:0] _GEN_294 = addr == 12'h301 ? pmpaddr0 : _GEN_273; // @[SIMD_CSR.scala 608:25 697:30]
  wire [63:0] _GEN_295 = addr == 12'h301 ? pmpaddr1 : _GEN_274; // @[SIMD_CSR.scala 609:25 697:30]
  wire [63:0] _GEN_296 = addr == 12'h301 ? pmpaddr2 : _GEN_275; // @[SIMD_CSR.scala 610:25 697:30]
  wire [63:0] _GEN_297 = addr == 12'h301 ? pmpaddr3 : _GEN_276; // @[SIMD_CSR.scala 611:25 697:30]
  wire [63:0] _GEN_298 = addr == 12'h301 ? vxsat : _GEN_277; // @[SIMD_CSR.scala 613:22 697:30]
  wire [63:0] _GEN_299 = addr == 12'h301 ? mipReg : _GEN_278; // @[SIMD_CSR.scala 583:24 697:30]
  wire  _GEN_300 = addr == 12'h301 ? 1'h0 : _GEN_279; // @[SIMD_CSR.scala 697:30]
  wire [63:0] _GEN_302 = addr == 12'h300 ? _GEN_12 : mstatus; // @[SIMD_CSR.scala 598:24 693:33]
  wire [63:0] _GEN_303 = addr == 12'h300 ? medeleg : _GEN_281; // @[SIMD_CSR.scala 600:24 693:33]
  wire [63:0] _GEN_304 = addr == 12'h300 ? mideleg : _GEN_282; // @[SIMD_CSR.scala 601:24 693:33]
  wire [63:0] _GEN_305 = addr == 12'h300 ? mie : _GEN_283; // @[SIMD_CSR.scala 581:20 693:33]
  wire [63:0] _GEN_306 = addr == 12'h300 ? mtvec : _GEN_284; // @[SIMD_CSR.scala 575:22 693:33]
  wire [63:0] _GEN_307 = addr == 12'h300 ? mcounteren : _GEN_285; // @[SIMD_CSR.scala 576:27 693:33]
  wire [63:0] _GEN_308 = addr == 12'h300 ? mscratch : _GEN_286; // @[SIMD_CSR.scala 602:25 693:33]
  wire [63:0] _GEN_309 = addr == 12'h300 ? mepc : _GEN_287; // @[SIMD_CSR.scala 579:17 693:33]
  wire [63:0] _GEN_310 = addr == 12'h300 ? mcause : _GEN_288; // @[SIMD_CSR.scala 577:23 693:33]
  wire [63:0] _GEN_311 = addr == 12'h300 ? mtval : _GEN_289; // @[SIMD_CSR.scala 578:22 693:33]
  wire [63:0] _GEN_312 = addr == 12'h300 ? pmpcfg0 : _GEN_290; // @[SIMD_CSR.scala 604:24 693:33]
  wire [63:0] _GEN_313 = addr == 12'h300 ? pmpcfg1 : _GEN_291; // @[SIMD_CSR.scala 605:24 693:33]
  wire [63:0] _GEN_314 = addr == 12'h300 ? pmpcfg2 : _GEN_292; // @[SIMD_CSR.scala 606:24 693:33]
  wire [63:0] _GEN_315 = addr == 12'h300 ? pmpcfg3 : _GEN_293; // @[SIMD_CSR.scala 607:24 693:33]
  wire [63:0] _GEN_316 = addr == 12'h300 ? pmpaddr0 : _GEN_294; // @[SIMD_CSR.scala 608:25 693:33]
  wire [63:0] _GEN_317 = addr == 12'h300 ? pmpaddr1 : _GEN_295; // @[SIMD_CSR.scala 609:25 693:33]
  wire [63:0] _GEN_318 = addr == 12'h300 ? pmpaddr2 : _GEN_296; // @[SIMD_CSR.scala 610:25 693:33]
  wire [63:0] _GEN_319 = addr == 12'h300 ? pmpaddr3 : _GEN_297; // @[SIMD_CSR.scala 611:25 693:33]
  wire [63:0] _GEN_320 = addr == 12'h300 ? vxsat : _GEN_298; // @[SIMD_CSR.scala 613:22 693:33]
  wire [63:0] _GEN_321 = addr == 12'h300 ? mipReg : _GEN_299; // @[SIMD_CSR.scala 583:24 693:33]
  wire  _GEN_322 = addr == 12'h300 ? 1'h0 : _GEN_300; // @[SIMD_CSR.scala 693:33]
  wire [63:0] _GEN_324 = addr == 12'h180 ? _GEN_10 : satp; // @[SIMD_CSR.scala 623:21 687:30]
  wire  _GEN_325 = addr == 12'h180 & _T_126; // @[SIMD_CSR.scala 687:30]
  wire [63:0] _GEN_326 = addr == 12'h180 ? mstatus : _GEN_302; // @[SIMD_CSR.scala 598:24 687:30]
  wire [63:0] _GEN_327 = addr == 12'h180 ? medeleg : _GEN_303; // @[SIMD_CSR.scala 600:24 687:30]
  wire [63:0] _GEN_328 = addr == 12'h180 ? mideleg : _GEN_304; // @[SIMD_CSR.scala 601:24 687:30]
  wire [63:0] _GEN_329 = addr == 12'h180 ? mie : _GEN_305; // @[SIMD_CSR.scala 581:20 687:30]
  wire [63:0] _GEN_330 = addr == 12'h180 ? mtvec : _GEN_306; // @[SIMD_CSR.scala 575:22 687:30]
  wire [63:0] _GEN_331 = addr == 12'h180 ? mcounteren : _GEN_307; // @[SIMD_CSR.scala 576:27 687:30]
  wire [63:0] _GEN_332 = addr == 12'h180 ? mscratch : _GEN_308; // @[SIMD_CSR.scala 602:25 687:30]
  wire [63:0] _GEN_333 = addr == 12'h180 ? mepc : _GEN_309; // @[SIMD_CSR.scala 579:17 687:30]
  wire [63:0] _GEN_334 = addr == 12'h180 ? mcause : _GEN_310; // @[SIMD_CSR.scala 577:23 687:30]
  wire [63:0] _GEN_335 = addr == 12'h180 ? mtval : _GEN_311; // @[SIMD_CSR.scala 578:22 687:30]
  wire [63:0] _GEN_336 = addr == 12'h180 ? pmpcfg0 : _GEN_312; // @[SIMD_CSR.scala 604:24 687:30]
  wire [63:0] _GEN_337 = addr == 12'h180 ? pmpcfg1 : _GEN_313; // @[SIMD_CSR.scala 605:24 687:30]
  wire [63:0] _GEN_338 = addr == 12'h180 ? pmpcfg2 : _GEN_314; // @[SIMD_CSR.scala 606:24 687:30]
  wire [63:0] _GEN_339 = addr == 12'h180 ? pmpcfg3 : _GEN_315; // @[SIMD_CSR.scala 607:24 687:30]
  wire [63:0] _GEN_340 = addr == 12'h180 ? pmpaddr0 : _GEN_316; // @[SIMD_CSR.scala 608:25 687:30]
  wire [63:0] _GEN_341 = addr == 12'h180 ? pmpaddr1 : _GEN_317; // @[SIMD_CSR.scala 609:25 687:30]
  wire [63:0] _GEN_342 = addr == 12'h180 ? pmpaddr2 : _GEN_318; // @[SIMD_CSR.scala 610:25 687:30]
  wire [63:0] _GEN_343 = addr == 12'h180 ? pmpaddr3 : _GEN_319; // @[SIMD_CSR.scala 611:25 687:30]
  wire [63:0] _GEN_344 = addr == 12'h180 ? vxsat : _GEN_320; // @[SIMD_CSR.scala 613:22 687:30]
  wire [63:0] _GEN_345 = addr == 12'h180 ? mipReg : _GEN_321; // @[SIMD_CSR.scala 583:24 687:30]
  wire  _GEN_346 = addr == 12'h180 ? 1'h0 : _GEN_322; // @[SIMD_CSR.scala 687:30]
  wire [63:0] _GEN_348 = addr == 12'h143 ? _GEN_9 : stval; // @[SIMD_CSR.scala 626:18 684:31]
  wire [63:0] _GEN_349 = addr == 12'h143 ? satp : _GEN_324; // @[SIMD_CSR.scala 623:21 684:31]
  wire  _GEN_350 = addr == 12'h143 ? 1'h0 : _GEN_325; // @[SIMD_CSR.scala 684:31]
  wire [63:0] _GEN_351 = addr == 12'h143 ? mstatus : _GEN_326; // @[SIMD_CSR.scala 598:24 684:31]
  wire [63:0] _GEN_352 = addr == 12'h143 ? medeleg : _GEN_327; // @[SIMD_CSR.scala 600:24 684:31]
  wire [63:0] _GEN_353 = addr == 12'h143 ? mideleg : _GEN_328; // @[SIMD_CSR.scala 601:24 684:31]
  wire [63:0] _GEN_354 = addr == 12'h143 ? mie : _GEN_329; // @[SIMD_CSR.scala 581:20 684:31]
  wire [63:0] _GEN_355 = addr == 12'h143 ? mtvec : _GEN_330; // @[SIMD_CSR.scala 575:22 684:31]
  wire [63:0] _GEN_356 = addr == 12'h143 ? mcounteren : _GEN_331; // @[SIMD_CSR.scala 576:27 684:31]
  wire [63:0] _GEN_357 = addr == 12'h143 ? mscratch : _GEN_332; // @[SIMD_CSR.scala 602:25 684:31]
  wire [63:0] _GEN_358 = addr == 12'h143 ? mepc : _GEN_333; // @[SIMD_CSR.scala 579:17 684:31]
  wire [63:0] _GEN_359 = addr == 12'h143 ? mcause : _GEN_334; // @[SIMD_CSR.scala 577:23 684:31]
  wire [63:0] _GEN_360 = addr == 12'h143 ? mtval : _GEN_335; // @[SIMD_CSR.scala 578:22 684:31]
  wire [63:0] _GEN_361 = addr == 12'h143 ? pmpcfg0 : _GEN_336; // @[SIMD_CSR.scala 604:24 684:31]
  wire [63:0] _GEN_362 = addr == 12'h143 ? pmpcfg1 : _GEN_337; // @[SIMD_CSR.scala 605:24 684:31]
  wire [63:0] _GEN_363 = addr == 12'h143 ? pmpcfg2 : _GEN_338; // @[SIMD_CSR.scala 606:24 684:31]
  wire [63:0] _GEN_364 = addr == 12'h143 ? pmpcfg3 : _GEN_339; // @[SIMD_CSR.scala 607:24 684:31]
  wire [63:0] _GEN_365 = addr == 12'h143 ? pmpaddr0 : _GEN_340; // @[SIMD_CSR.scala 608:25 684:31]
  wire [63:0] _GEN_366 = addr == 12'h143 ? pmpaddr1 : _GEN_341; // @[SIMD_CSR.scala 609:25 684:31]
  wire [63:0] _GEN_367 = addr == 12'h143 ? pmpaddr2 : _GEN_342; // @[SIMD_CSR.scala 610:25 684:31]
  wire [63:0] _GEN_368 = addr == 12'h143 ? pmpaddr3 : _GEN_343; // @[SIMD_CSR.scala 611:25 684:31]
  wire [63:0] _GEN_369 = addr == 12'h143 ? vxsat : _GEN_344; // @[SIMD_CSR.scala 613:22 684:31]
  wire [63:0] _GEN_370 = addr == 12'h143 ? mipReg : _GEN_345; // @[SIMD_CSR.scala 583:24 684:31]
  wire  _GEN_371 = addr == 12'h143 ? 1'h0 : _GEN_346; // @[SIMD_CSR.scala 684:31]
  wire [63:0] _GEN_373 = addr == 12'h142 ? _GEN_8 : scause; // @[SIMD_CSR.scala 625:23 681:32]
  wire [63:0] _GEN_374 = addr == 12'h142 ? stval : _GEN_348; // @[SIMD_CSR.scala 626:18 681:32]
  wire [63:0] _GEN_375 = addr == 12'h142 ? satp : _GEN_349; // @[SIMD_CSR.scala 623:21 681:32]
  wire  _GEN_376 = addr == 12'h142 ? 1'h0 : _GEN_350; // @[SIMD_CSR.scala 681:32]
  wire [63:0] _GEN_377 = addr == 12'h142 ? mstatus : _GEN_351; // @[SIMD_CSR.scala 598:24 681:32]
  wire [63:0] _GEN_378 = addr == 12'h142 ? medeleg : _GEN_352; // @[SIMD_CSR.scala 600:24 681:32]
  wire [63:0] _GEN_379 = addr == 12'h142 ? mideleg : _GEN_353; // @[SIMD_CSR.scala 601:24 681:32]
  wire [63:0] _GEN_380 = addr == 12'h142 ? mie : _GEN_354; // @[SIMD_CSR.scala 581:20 681:32]
  wire [63:0] _GEN_381 = addr == 12'h142 ? mtvec : _GEN_355; // @[SIMD_CSR.scala 575:22 681:32]
  wire [63:0] _GEN_382 = addr == 12'h142 ? mcounteren : _GEN_356; // @[SIMD_CSR.scala 576:27 681:32]
  wire [63:0] _GEN_383 = addr == 12'h142 ? mscratch : _GEN_357; // @[SIMD_CSR.scala 602:25 681:32]
  wire [63:0] _GEN_384 = addr == 12'h142 ? mepc : _GEN_358; // @[SIMD_CSR.scala 579:17 681:32]
  wire [63:0] _GEN_385 = addr == 12'h142 ? mcause : _GEN_359; // @[SIMD_CSR.scala 577:23 681:32]
  wire [63:0] _GEN_386 = addr == 12'h142 ? mtval : _GEN_360; // @[SIMD_CSR.scala 578:22 681:32]
  wire [63:0] _GEN_387 = addr == 12'h142 ? pmpcfg0 : _GEN_361; // @[SIMD_CSR.scala 604:24 681:32]
  wire [63:0] _GEN_388 = addr == 12'h142 ? pmpcfg1 : _GEN_362; // @[SIMD_CSR.scala 605:24 681:32]
  wire [63:0] _GEN_389 = addr == 12'h142 ? pmpcfg2 : _GEN_363; // @[SIMD_CSR.scala 606:24 681:32]
  wire [63:0] _GEN_390 = addr == 12'h142 ? pmpcfg3 : _GEN_364; // @[SIMD_CSR.scala 607:24 681:32]
  wire [63:0] _GEN_391 = addr == 12'h142 ? pmpaddr0 : _GEN_365; // @[SIMD_CSR.scala 608:25 681:32]
  wire [63:0] _GEN_392 = addr == 12'h142 ? pmpaddr1 : _GEN_366; // @[SIMD_CSR.scala 609:25 681:32]
  wire [63:0] _GEN_393 = addr == 12'h142 ? pmpaddr2 : _GEN_367; // @[SIMD_CSR.scala 610:25 681:32]
  wire [63:0] _GEN_394 = addr == 12'h142 ? pmpaddr3 : _GEN_368; // @[SIMD_CSR.scala 611:25 681:32]
  wire [63:0] _GEN_395 = addr == 12'h142 ? vxsat : _GEN_369; // @[SIMD_CSR.scala 613:22 681:32]
  wire [63:0] _GEN_396 = addr == 12'h142 ? mipReg : _GEN_370; // @[SIMD_CSR.scala 583:24 681:32]
  wire  _GEN_397 = addr == 12'h142 ? 1'h0 : _GEN_371; // @[SIMD_CSR.scala 681:32]
  wire [63:0] _GEN_399 = addr == 12'h141 ? _GEN_7 : sepc; // @[SIMD_CSR.scala 624:21 678:30]
  wire [63:0] _GEN_400 = addr == 12'h141 ? scause : _GEN_373; // @[SIMD_CSR.scala 625:23 678:30]
  wire [63:0] _GEN_401 = addr == 12'h141 ? stval : _GEN_374; // @[SIMD_CSR.scala 626:18 678:30]
  wire [63:0] _GEN_402 = addr == 12'h141 ? satp : _GEN_375; // @[SIMD_CSR.scala 623:21 678:30]
  wire  _GEN_403 = addr == 12'h141 ? 1'h0 : _GEN_376; // @[SIMD_CSR.scala 678:30]
  wire [63:0] _GEN_404 = addr == 12'h141 ? mstatus : _GEN_377; // @[SIMD_CSR.scala 598:24 678:30]
  wire [63:0] _GEN_405 = addr == 12'h141 ? medeleg : _GEN_378; // @[SIMD_CSR.scala 600:24 678:30]
  wire [63:0] _GEN_406 = addr == 12'h141 ? mideleg : _GEN_379; // @[SIMD_CSR.scala 601:24 678:30]
  wire [63:0] _GEN_407 = addr == 12'h141 ? mie : _GEN_380; // @[SIMD_CSR.scala 581:20 678:30]
  wire [63:0] _GEN_408 = addr == 12'h141 ? mtvec : _GEN_381; // @[SIMD_CSR.scala 575:22 678:30]
  wire [63:0] _GEN_409 = addr == 12'h141 ? mcounteren : _GEN_382; // @[SIMD_CSR.scala 576:27 678:30]
  wire [63:0] _GEN_410 = addr == 12'h141 ? mscratch : _GEN_383; // @[SIMD_CSR.scala 602:25 678:30]
  wire [63:0] _GEN_411 = addr == 12'h141 ? mepc : _GEN_384; // @[SIMD_CSR.scala 579:17 678:30]
  wire [63:0] _GEN_412 = addr == 12'h141 ? mcause : _GEN_385; // @[SIMD_CSR.scala 577:23 678:30]
  wire [63:0] _GEN_413 = addr == 12'h141 ? mtval : _GEN_386; // @[SIMD_CSR.scala 578:22 678:30]
  wire [63:0] _GEN_414 = addr == 12'h141 ? pmpcfg0 : _GEN_387; // @[SIMD_CSR.scala 604:24 678:30]
  wire [63:0] _GEN_415 = addr == 12'h141 ? pmpcfg1 : _GEN_388; // @[SIMD_CSR.scala 605:24 678:30]
  wire [63:0] _GEN_416 = addr == 12'h141 ? pmpcfg2 : _GEN_389; // @[SIMD_CSR.scala 606:24 678:30]
  wire [63:0] _GEN_417 = addr == 12'h141 ? pmpcfg3 : _GEN_390; // @[SIMD_CSR.scala 607:24 678:30]
  wire [63:0] _GEN_418 = addr == 12'h141 ? pmpaddr0 : _GEN_391; // @[SIMD_CSR.scala 608:25 678:30]
  wire [63:0] _GEN_419 = addr == 12'h141 ? pmpaddr1 : _GEN_392; // @[SIMD_CSR.scala 609:25 678:30]
  wire [63:0] _GEN_420 = addr == 12'h141 ? pmpaddr2 : _GEN_393; // @[SIMD_CSR.scala 610:25 678:30]
  wire [63:0] _GEN_421 = addr == 12'h141 ? pmpaddr3 : _GEN_394; // @[SIMD_CSR.scala 611:25 678:30]
  wire [63:0] _GEN_422 = addr == 12'h141 ? vxsat : _GEN_395; // @[SIMD_CSR.scala 613:22 678:30]
  wire [63:0] _GEN_423 = addr == 12'h141 ? mipReg : _GEN_396; // @[SIMD_CSR.scala 583:24 678:30]
  wire  _GEN_424 = addr == 12'h141 ? 1'h0 : _GEN_397; // @[SIMD_CSR.scala 678:30]
  wire [63:0] _GEN_426 = addr == 12'h140 ? _GEN_6 : sscratch; // @[SIMD_CSR.scala 627:25 675:34]
  wire [63:0] _GEN_427 = addr == 12'h140 ? sepc : _GEN_399; // @[SIMD_CSR.scala 624:21 675:34]
  wire [63:0] _GEN_428 = addr == 12'h140 ? scause : _GEN_400; // @[SIMD_CSR.scala 625:23 675:34]
  wire [63:0] _GEN_429 = addr == 12'h140 ? stval : _GEN_401; // @[SIMD_CSR.scala 626:18 675:34]
  wire [63:0] _GEN_430 = addr == 12'h140 ? satp : _GEN_402; // @[SIMD_CSR.scala 623:21 675:34]
  wire  _GEN_431 = addr == 12'h140 ? 1'h0 : _GEN_403; // @[SIMD_CSR.scala 675:34]
  wire [63:0] _GEN_432 = addr == 12'h140 ? mstatus : _GEN_404; // @[SIMD_CSR.scala 598:24 675:34]
  wire [63:0] _GEN_433 = addr == 12'h140 ? medeleg : _GEN_405; // @[SIMD_CSR.scala 600:24 675:34]
  wire [63:0] _GEN_434 = addr == 12'h140 ? mideleg : _GEN_406; // @[SIMD_CSR.scala 601:24 675:34]
  wire [63:0] _GEN_435 = addr == 12'h140 ? mie : _GEN_407; // @[SIMD_CSR.scala 581:20 675:34]
  wire [63:0] _GEN_436 = addr == 12'h140 ? mtvec : _GEN_408; // @[SIMD_CSR.scala 575:22 675:34]
  wire [63:0] _GEN_437 = addr == 12'h140 ? mcounteren : _GEN_409; // @[SIMD_CSR.scala 576:27 675:34]
  wire [63:0] _GEN_438 = addr == 12'h140 ? mscratch : _GEN_410; // @[SIMD_CSR.scala 602:25 675:34]
  wire [63:0] _GEN_439 = addr == 12'h140 ? mepc : _GEN_411; // @[SIMD_CSR.scala 579:17 675:34]
  wire [63:0] _GEN_440 = addr == 12'h140 ? mcause : _GEN_412; // @[SIMD_CSR.scala 577:23 675:34]
  wire [63:0] _GEN_441 = addr == 12'h140 ? mtval : _GEN_413; // @[SIMD_CSR.scala 578:22 675:34]
  wire [63:0] _GEN_442 = addr == 12'h140 ? pmpcfg0 : _GEN_414; // @[SIMD_CSR.scala 604:24 675:34]
  wire [63:0] _GEN_443 = addr == 12'h140 ? pmpcfg1 : _GEN_415; // @[SIMD_CSR.scala 605:24 675:34]
  wire [63:0] _GEN_444 = addr == 12'h140 ? pmpcfg2 : _GEN_416; // @[SIMD_CSR.scala 606:24 675:34]
  wire [63:0] _GEN_445 = addr == 12'h140 ? pmpcfg3 : _GEN_417; // @[SIMD_CSR.scala 607:24 675:34]
  wire [63:0] _GEN_446 = addr == 12'h140 ? pmpaddr0 : _GEN_418; // @[SIMD_CSR.scala 608:25 675:34]
  wire [63:0] _GEN_447 = addr == 12'h140 ? pmpaddr1 : _GEN_419; // @[SIMD_CSR.scala 609:25 675:34]
  wire [63:0] _GEN_448 = addr == 12'h140 ? pmpaddr2 : _GEN_420; // @[SIMD_CSR.scala 610:25 675:34]
  wire [63:0] _GEN_449 = addr == 12'h140 ? pmpaddr3 : _GEN_421; // @[SIMD_CSR.scala 611:25 675:34]
  wire [63:0] _GEN_450 = addr == 12'h140 ? vxsat : _GEN_422; // @[SIMD_CSR.scala 613:22 675:34]
  wire [63:0] _GEN_451 = addr == 12'h140 ? mipReg : _GEN_423; // @[SIMD_CSR.scala 583:24 675:34]
  wire  _GEN_452 = addr == 12'h140 ? 1'h0 : _GEN_424; // @[SIMD_CSR.scala 675:34]
  wire [63:0] _GEN_454 = addr == 12'h106 ? _GEN_5 : scounteren; // @[SIMD_CSR.scala 628:27 672:36]
  wire [63:0] _GEN_455 = addr == 12'h106 ? sscratch : _GEN_426; // @[SIMD_CSR.scala 627:25 672:36]
  wire [63:0] _GEN_456 = addr == 12'h106 ? sepc : _GEN_427; // @[SIMD_CSR.scala 624:21 672:36]
  wire [63:0] _GEN_457 = addr == 12'h106 ? scause : _GEN_428; // @[SIMD_CSR.scala 625:23 672:36]
  wire [63:0] _GEN_458 = addr == 12'h106 ? stval : _GEN_429; // @[SIMD_CSR.scala 626:18 672:36]
  wire [63:0] _GEN_459 = addr == 12'h106 ? satp : _GEN_430; // @[SIMD_CSR.scala 623:21 672:36]
  wire  _GEN_460 = addr == 12'h106 ? 1'h0 : _GEN_431; // @[SIMD_CSR.scala 672:36]
  wire [63:0] _GEN_461 = addr == 12'h106 ? mstatus : _GEN_432; // @[SIMD_CSR.scala 598:24 672:36]
  wire [63:0] _GEN_462 = addr == 12'h106 ? medeleg : _GEN_433; // @[SIMD_CSR.scala 600:24 672:36]
  wire [63:0] _GEN_463 = addr == 12'h106 ? mideleg : _GEN_434; // @[SIMD_CSR.scala 601:24 672:36]
  wire [63:0] _GEN_464 = addr == 12'h106 ? mie : _GEN_435; // @[SIMD_CSR.scala 581:20 672:36]
  wire [63:0] _GEN_465 = addr == 12'h106 ? mtvec : _GEN_436; // @[SIMD_CSR.scala 575:22 672:36]
  wire [63:0] _GEN_466 = addr == 12'h106 ? mcounteren : _GEN_437; // @[SIMD_CSR.scala 576:27 672:36]
  wire [63:0] _GEN_467 = addr == 12'h106 ? mscratch : _GEN_438; // @[SIMD_CSR.scala 602:25 672:36]
  wire [63:0] _GEN_468 = addr == 12'h106 ? mepc : _GEN_439; // @[SIMD_CSR.scala 579:17 672:36]
  wire [63:0] _GEN_469 = addr == 12'h106 ? mcause : _GEN_440; // @[SIMD_CSR.scala 577:23 672:36]
  wire [63:0] _GEN_470 = addr == 12'h106 ? mtval : _GEN_441; // @[SIMD_CSR.scala 578:22 672:36]
  wire [63:0] _GEN_471 = addr == 12'h106 ? pmpcfg0 : _GEN_442; // @[SIMD_CSR.scala 604:24 672:36]
  wire [63:0] _GEN_472 = addr == 12'h106 ? pmpcfg1 : _GEN_443; // @[SIMD_CSR.scala 605:24 672:36]
  wire [63:0] _GEN_473 = addr == 12'h106 ? pmpcfg2 : _GEN_444; // @[SIMD_CSR.scala 606:24 672:36]
  wire [63:0] _GEN_474 = addr == 12'h106 ? pmpcfg3 : _GEN_445; // @[SIMD_CSR.scala 607:24 672:36]
  wire [63:0] _GEN_475 = addr == 12'h106 ? pmpaddr0 : _GEN_446; // @[SIMD_CSR.scala 608:25 672:36]
  wire [63:0] _GEN_476 = addr == 12'h106 ? pmpaddr1 : _GEN_447; // @[SIMD_CSR.scala 609:25 672:36]
  wire [63:0] _GEN_477 = addr == 12'h106 ? pmpaddr2 : _GEN_448; // @[SIMD_CSR.scala 610:25 672:36]
  wire [63:0] _GEN_478 = addr == 12'h106 ? pmpaddr3 : _GEN_449; // @[SIMD_CSR.scala 611:25 672:36]
  wire [63:0] _GEN_479 = addr == 12'h106 ? vxsat : _GEN_450; // @[SIMD_CSR.scala 613:22 672:36]
  wire [63:0] _GEN_480 = addr == 12'h106 ? mipReg : _GEN_451; // @[SIMD_CSR.scala 583:24 672:36]
  wire  _GEN_481 = addr == 12'h106 ? 1'h0 : _GEN_452; // @[SIMD_CSR.scala 672:36]
  wire [63:0] _GEN_486 = addr == 12'h105 ? sepc : _GEN_456; // @[SIMD_CSR.scala 624:21 669:31]
  wire [63:0] _GEN_487 = addr == 12'h105 ? scause : _GEN_457; // @[SIMD_CSR.scala 625:23 669:31]
  wire [63:0] _GEN_488 = addr == 12'h105 ? stval : _GEN_458; // @[SIMD_CSR.scala 626:18 669:31]
  wire  _GEN_490 = addr == 12'h105 ? 1'h0 : _GEN_460; // @[SIMD_CSR.scala 669:31]
  wire [63:0] _GEN_491 = addr == 12'h105 ? mstatus : _GEN_461; // @[SIMD_CSR.scala 598:24 669:31]
  wire [63:0] _GEN_498 = addr == 12'h105 ? mepc : _GEN_468; // @[SIMD_CSR.scala 579:17 669:31]
  wire [63:0] _GEN_499 = addr == 12'h105 ? mcause : _GEN_469; // @[SIMD_CSR.scala 577:23 669:31]
  wire [63:0] _GEN_500 = addr == 12'h105 ? mtval : _GEN_470; // @[SIMD_CSR.scala 578:22 669:31]
  wire [63:0] _GEN_509 = addr == 12'h105 ? vxsat : _GEN_479; // @[SIMD_CSR.scala 613:22 669:31]
  wire  _GEN_511 = addr == 12'h105 ? 1'h0 : _GEN_481; // @[SIMD_CSR.scala 669:31]
  wire [63:0] _GEN_517 = addr == 12'h104 ? sepc : _GEN_486; // @[SIMD_CSR.scala 624:21 666:29]
  wire [63:0] _GEN_518 = addr == 12'h104 ? scause : _GEN_487; // @[SIMD_CSR.scala 625:23 666:29]
  wire [63:0] _GEN_519 = addr == 12'h104 ? stval : _GEN_488; // @[SIMD_CSR.scala 626:18 666:29]
  wire  _GEN_521 = addr == 12'h104 ? 1'h0 : _GEN_490; // @[SIMD_CSR.scala 666:29]
  wire [63:0] _GEN_522 = addr == 12'h104 ? mstatus : _GEN_491; // @[SIMD_CSR.scala 598:24 666:29]
  wire [63:0] _GEN_528 = addr == 12'h104 ? mepc : _GEN_498; // @[SIMD_CSR.scala 579:17 666:29]
  wire [63:0] _GEN_529 = addr == 12'h104 ? mcause : _GEN_499; // @[SIMD_CSR.scala 577:23 666:29]
  wire [63:0] _GEN_530 = addr == 12'h104 ? mtval : _GEN_500; // @[SIMD_CSR.scala 578:22 666:29]
  wire  _GEN_541 = addr == 12'h104 ? 1'h0 : _GEN_511; // @[SIMD_CSR.scala 666:29]
  wire [63:0] _GEN_548 = addr == 12'h100 ? sepc : _GEN_517; // @[SIMD_CSR.scala 624:21 662:27]
  wire [63:0] _GEN_549 = addr == 12'h100 ? scause : _GEN_518; // @[SIMD_CSR.scala 625:23 662:27]
  wire [63:0] _GEN_550 = addr == 12'h100 ? stval : _GEN_519; // @[SIMD_CSR.scala 626:18 662:27]
  wire  resetSatp = addr == 12'h100 ? 1'h0 : _GEN_521; // @[SIMD_CSR.scala 662:27]
  wire [63:0] _GEN_558 = addr == 12'h100 ? mepc : _GEN_528; // @[SIMD_CSR.scala 579:17 662:27]
  wire [63:0] _GEN_559 = addr == 12'h100 ? mcause : _GEN_529; // @[SIMD_CSR.scala 577:23 662:27]
  wire [63:0] _GEN_560 = addr == 12'h100 ? mtval : _GEN_530; // @[SIMD_CSR.scala 578:22 662:27]
  wire  isIllegalAddr = addr == 12'h100 ? 1'h0 : _GEN_541; // @[SIMD_CSR.scala 662:27]
  wire  isMret = _T_156 & JumpType; // @[SIMD_CSR.scala 778:35]
  wire  isSret = addr == 12'h102 & JumpType; // @[SIMD_CSR.scala 779:35]
  wire  isUret = addr == 12'h2 & JumpType; // @[SIMD_CSR.scala 780:35]
  wire  isIllegalSret = isSret & mstatusStruct_tsr; // @[SIMD_CSR.scala 781:30]
  wire  isRet = io_in_valid & _T_55 & (isMret | isSret | isUret) & ~isIllegalSret; // @[SIMD_CSR.scala 782:65]
  wire  _T_247 = priviledgeMode < 2'h3; // @[SIMD_CSR.scala 791:63]
  wire  _T_248 = priviledgeMode == 2'h1; // @[SIMD_CSR.scala 791:89]
  wire  _T_254 = ~mideleg[0] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_0 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_254; // @[SIMD_CSR.scala 791:47]
  wire  _T_263 = ~mideleg[1] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_1 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_263; // @[SIMD_CSR.scala 791:47]
  wire  _T_272 = ~mideleg[2] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_2 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_272; // @[SIMD_CSR.scala 791:47]
  wire  _T_281 = ~mideleg[3] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_3 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_281; // @[SIMD_CSR.scala 791:47]
  wire  _T_290 = ~mideleg[4] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_4 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_290; // @[SIMD_CSR.scala 791:47]
  wire  _T_299 = ~mideleg[5] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_5 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_299; // @[SIMD_CSR.scala 791:47]
  wire  _T_308 = ~mideleg[6] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_6 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_308; // @[SIMD_CSR.scala 791:47]
  wire  _T_317 = ~mideleg[7] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_7 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_317; // @[SIMD_CSR.scala 791:47]
  wire  _T_326 = ~mideleg[8] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_8 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_326; // @[SIMD_CSR.scala 791:47]
  wire  _T_335 = ~mideleg[9] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_9 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _T_335; // @[SIMD_CSR.scala 791:47]
  wire  _T_344 = ~mideleg[10] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_10 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1
     : _T_344; // @[SIMD_CSR.scala 791:47]
  wire  _T_353 = ~mideleg[11] & mstatusStruct_ie_m; // @[SIMD_CSR.scala 792:87]
  wire  intrVecEnable_11 = priviledgeMode < 2'h3 ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1
     : _T_353; // @[SIMD_CSR.scala 791:47]
  wire [63:0] _GEN_920 = {{52'd0}, mie[11:0]}; // @[SIMD_CSR.scala 794:27]
  wire [63:0] _T_357 = _GEN_920 & _T_209; // @[SIMD_CSR.scala 794:27]
  wire [5:0] lo_4 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,intrVecEnable_0}; // @[SIMD_CSR.scala 794:52]
  wire [11:0] _T_358 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,lo_4}; // @[SIMD_CSR.scala 794:52]
  wire [63:0] _GEN_921 = {{52'd0}, _T_358}; // @[SIMD_CSR.scala 794:36]
  wire [63:0] intrVec = _T_357 & _GEN_921; // @[SIMD_CSR.scala 794:36]
  wire [3:0] _T_359 = io_cfIn_intrVec_3 ? 4'h3 : 4'hb; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_574 = 4'h1 == _T_359 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_575 = 4'h2 == _T_359 ? io_cfIn_intrVec_2 : _GEN_574; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_576 = 4'h3 == _T_359 ? io_cfIn_intrVec_3 : _GEN_575; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_577 = 4'h4 == _T_359 ? io_cfIn_intrVec_4 : _GEN_576; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_578 = 4'h5 == _T_359 ? io_cfIn_intrVec_5 : _GEN_577; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_579 = 4'h6 == _T_359 ? io_cfIn_intrVec_6 : _GEN_578; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_580 = 4'h7 == _T_359 ? io_cfIn_intrVec_7 : _GEN_579; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_581 = 4'h8 == _T_359 ? io_cfIn_intrVec_8 : _GEN_580; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_582 = 4'h9 == _T_359 ? io_cfIn_intrVec_9 : _GEN_581; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_583 = 4'ha == _T_359 ? io_cfIn_intrVec_10 : _GEN_582; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_584 = 4'hb == _T_359 ? io_cfIn_intrVec_11 : _GEN_583; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] _T_360 = _GEN_584 ? _T_359 : 4'h7; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_586 = 4'h1 == _T_360 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_587 = 4'h2 == _T_360 ? io_cfIn_intrVec_2 : _GEN_586; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_588 = 4'h3 == _T_360 ? io_cfIn_intrVec_3 : _GEN_587; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_589 = 4'h4 == _T_360 ? io_cfIn_intrVec_4 : _GEN_588; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_590 = 4'h5 == _T_360 ? io_cfIn_intrVec_5 : _GEN_589; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_591 = 4'h6 == _T_360 ? io_cfIn_intrVec_6 : _GEN_590; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_592 = 4'h7 == _T_360 ? io_cfIn_intrVec_7 : _GEN_591; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_593 = 4'h8 == _T_360 ? io_cfIn_intrVec_8 : _GEN_592; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_594 = 4'h9 == _T_360 ? io_cfIn_intrVec_9 : _GEN_593; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_595 = 4'ha == _T_360 ? io_cfIn_intrVec_10 : _GEN_594; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_596 = 4'hb == _T_360 ? io_cfIn_intrVec_11 : _GEN_595; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] _T_361 = _GEN_596 ? _T_360 : 4'h1; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_598 = 4'h1 == _T_361 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_599 = 4'h2 == _T_361 ? io_cfIn_intrVec_2 : _GEN_598; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_600 = 4'h3 == _T_361 ? io_cfIn_intrVec_3 : _GEN_599; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_601 = 4'h4 == _T_361 ? io_cfIn_intrVec_4 : _GEN_600; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_602 = 4'h5 == _T_361 ? io_cfIn_intrVec_5 : _GEN_601; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_603 = 4'h6 == _T_361 ? io_cfIn_intrVec_6 : _GEN_602; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_604 = 4'h7 == _T_361 ? io_cfIn_intrVec_7 : _GEN_603; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_605 = 4'h8 == _T_361 ? io_cfIn_intrVec_8 : _GEN_604; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_606 = 4'h9 == _T_361 ? io_cfIn_intrVec_9 : _GEN_605; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_607 = 4'ha == _T_361 ? io_cfIn_intrVec_10 : _GEN_606; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_608 = 4'hb == _T_361 ? io_cfIn_intrVec_11 : _GEN_607; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] _T_362 = _GEN_608 ? _T_361 : 4'h9; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_610 = 4'h1 == _T_362 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_611 = 4'h2 == _T_362 ? io_cfIn_intrVec_2 : _GEN_610; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_612 = 4'h3 == _T_362 ? io_cfIn_intrVec_3 : _GEN_611; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_613 = 4'h4 == _T_362 ? io_cfIn_intrVec_4 : _GEN_612; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_614 = 4'h5 == _T_362 ? io_cfIn_intrVec_5 : _GEN_613; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_615 = 4'h6 == _T_362 ? io_cfIn_intrVec_6 : _GEN_614; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_616 = 4'h7 == _T_362 ? io_cfIn_intrVec_7 : _GEN_615; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_617 = 4'h8 == _T_362 ? io_cfIn_intrVec_8 : _GEN_616; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_618 = 4'h9 == _T_362 ? io_cfIn_intrVec_9 : _GEN_617; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_619 = 4'ha == _T_362 ? io_cfIn_intrVec_10 : _GEN_618; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_620 = 4'hb == _T_362 ? io_cfIn_intrVec_11 : _GEN_619; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] _T_363 = _GEN_620 ? _T_362 : 4'h5; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_622 = 4'h1 == _T_363 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_623 = 4'h2 == _T_363 ? io_cfIn_intrVec_2 : _GEN_622; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_624 = 4'h3 == _T_363 ? io_cfIn_intrVec_3 : _GEN_623; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_625 = 4'h4 == _T_363 ? io_cfIn_intrVec_4 : _GEN_624; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_626 = 4'h5 == _T_363 ? io_cfIn_intrVec_5 : _GEN_625; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_627 = 4'h6 == _T_363 ? io_cfIn_intrVec_6 : _GEN_626; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_628 = 4'h7 == _T_363 ? io_cfIn_intrVec_7 : _GEN_627; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_629 = 4'h8 == _T_363 ? io_cfIn_intrVec_8 : _GEN_628; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_630 = 4'h9 == _T_363 ? io_cfIn_intrVec_9 : _GEN_629; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_631 = 4'ha == _T_363 ? io_cfIn_intrVec_10 : _GEN_630; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_632 = 4'hb == _T_363 ? io_cfIn_intrVec_11 : _GEN_631; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] _T_364 = _GEN_632 ? _T_363 : 4'h0; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_634 = 4'h1 == _T_364 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_635 = 4'h2 == _T_364 ? io_cfIn_intrVec_2 : _GEN_634; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_636 = 4'h3 == _T_364 ? io_cfIn_intrVec_3 : _GEN_635; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_637 = 4'h4 == _T_364 ? io_cfIn_intrVec_4 : _GEN_636; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_638 = 4'h5 == _T_364 ? io_cfIn_intrVec_5 : _GEN_637; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_639 = 4'h6 == _T_364 ? io_cfIn_intrVec_6 : _GEN_638; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_640 = 4'h7 == _T_364 ? io_cfIn_intrVec_7 : _GEN_639; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_641 = 4'h8 == _T_364 ? io_cfIn_intrVec_8 : _GEN_640; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_642 = 4'h9 == _T_364 ? io_cfIn_intrVec_9 : _GEN_641; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_643 = 4'ha == _T_364 ? io_cfIn_intrVec_10 : _GEN_642; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_644 = 4'hb == _T_364 ? io_cfIn_intrVec_11 : _GEN_643; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] _T_365 = _GEN_644 ? _T_364 : 4'h8; // @[SIMD_CSR.scala 795:63]
  wire  _GEN_646 = 4'h1 == _T_365 ? io_cfIn_intrVec_1 : io_cfIn_intrVec_0; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_647 = 4'h2 == _T_365 ? io_cfIn_intrVec_2 : _GEN_646; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_648 = 4'h3 == _T_365 ? io_cfIn_intrVec_3 : _GEN_647; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_649 = 4'h4 == _T_365 ? io_cfIn_intrVec_4 : _GEN_648; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_650 = 4'h5 == _T_365 ? io_cfIn_intrVec_5 : _GEN_649; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_651 = 4'h6 == _T_365 ? io_cfIn_intrVec_6 : _GEN_650; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_652 = 4'h7 == _T_365 ? io_cfIn_intrVec_7 : _GEN_651; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_653 = 4'h8 == _T_365 ? io_cfIn_intrVec_8 : _GEN_652; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_654 = 4'h9 == _T_365 ? io_cfIn_intrVec_9 : _GEN_653; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_655 = 4'ha == _T_365 ? io_cfIn_intrVec_10 : _GEN_654; // @[SIMD_CSR.scala 795:{63,63}]
  wire  _GEN_656 = 4'hb == _T_365 ? io_cfIn_intrVec_11 : _GEN_655; // @[SIMD_CSR.scala 795:{63,63}]
  wire [3:0] intrNO = _GEN_656 ? _T_365 : 4'h4; // @[SIMD_CSR.scala 795:63]
  wire [5:0] lo_5 = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,
    io_cfIn_intrVec_0}; // @[SIMD_CSR.scala 796:35]
  wire [11:0] _T_366 = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,io_cfIn_intrVec_7,
    io_cfIn_intrVec_6,lo_5}; // @[SIMD_CSR.scala 796:35]
  wire  raiseIntr = |_T_366; // @[SIMD_CSR.scala 796:42]
  wire  csrExceptionVec_3 = io_in_valid & addr == 12'h1 & JumpType; // @[SIMD_CSR.scala 801:69]
  wire  _T_380 = addr == 12'h0; // @[SIMD_CSR.scala 802:78]
  wire  csrExceptionVec_11 = priviledgeMode == 2'h3 & io_in_valid & addr == 12'h0 & JumpType; // @[SIMD_CSR.scala 802:92]
  wire  csrExceptionVec_9 = _T_248 & io_in_valid & _T_380 & JumpType; // @[SIMD_CSR.scala 803:92]
  wire  csrExceptionVec_8 = priviledgeMode == 2'h0 & io_in_valid & _T_380 & JumpType; // @[SIMD_CSR.scala 804:92]
  wire  csrExceptionVec_2 = isIllegalAddr | isIllegalWrite | isIllegalMode | isIllegalSret | io_cfIn_exceptionVec_2; // @[SIMD_CSR.scala 805:102]
  wire  csrExceptionVec_13 = io_dmemMMU_loadPF | io_cfIn_exceptionVec_13; // @[SIMD_CSR.scala 806:55]
  wire  csrExceptionVec_15 = io_dmemMMU_storePF | io_cfIn_exceptionVec_15; // @[SIMD_CSR.scala 807:57]
  wire [7:0] lo_7 = {1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,csrExceptionVec_3,csrExceptionVec_2,
    io_cfIn_exceptionVec_1,1'h0}; // @[SIMD_CSR.scala 808:40]
  wire [15:0] _T_399 = {csrExceptionVec_15,1'h0,csrExceptionVec_13,io_cfIn_exceptionVec_12,csrExceptionVec_11,1'h0,
    csrExceptionVec_9,csrExceptionVec_8,lo_7}; // @[SIMD_CSR.scala 808:40]
  wire  raiseException = |_T_399; // @[SIMD_CSR.scala 808:47]
  wire [3:0] _T_400 = csrExceptionVec_3 ? 4'h3 : 4'hc; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_659 = 4'h2 == _T_400 ? csrExceptionVec_2 : 4'h1 == _T_400 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_660 = 4'h3 == _T_400 ? csrExceptionVec_3 : _GEN_659; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_661 = 4'h4 == _T_400 ? io_cfIn_exceptionVec_4 : _GEN_660; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_662 = 4'h5 == _T_400 ? 1'h0 : _GEN_661; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_663 = 4'h6 == _T_400 ? io_cfIn_exceptionVec_6 : _GEN_662; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_664 = 4'h7 == _T_400 ? 1'h0 : _GEN_663; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_665 = 4'h8 == _T_400 ? csrExceptionVec_8 : _GEN_664; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_666 = 4'h9 == _T_400 ? csrExceptionVec_9 : _GEN_665; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_667 = 4'ha == _T_400 ? 1'h0 : _GEN_666; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_668 = 4'hb == _T_400 ? csrExceptionVec_11 : _GEN_667; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_669 = 4'hc == _T_400 ? io_cfIn_exceptionVec_12 : _GEN_668; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_670 = 4'hd == _T_400 ? csrExceptionVec_13 : _GEN_669; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_671 = 4'he == _T_400 ? 1'h0 : _GEN_670; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_672 = 4'hf == _T_400 ? csrExceptionVec_15 : _GEN_671; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_401 = _GEN_672 ? _T_400 : 4'h1; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_675 = 4'h2 == _T_401 ? csrExceptionVec_2 : 4'h1 == _T_401 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_676 = 4'h3 == _T_401 ? csrExceptionVec_3 : _GEN_675; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_677 = 4'h4 == _T_401 ? io_cfIn_exceptionVec_4 : _GEN_676; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_678 = 4'h5 == _T_401 ? 1'h0 : _GEN_677; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_679 = 4'h6 == _T_401 ? io_cfIn_exceptionVec_6 : _GEN_678; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_680 = 4'h7 == _T_401 ? 1'h0 : _GEN_679; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_681 = 4'h8 == _T_401 ? csrExceptionVec_8 : _GEN_680; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_682 = 4'h9 == _T_401 ? csrExceptionVec_9 : _GEN_681; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_683 = 4'ha == _T_401 ? 1'h0 : _GEN_682; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_684 = 4'hb == _T_401 ? csrExceptionVec_11 : _GEN_683; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_685 = 4'hc == _T_401 ? io_cfIn_exceptionVec_12 : _GEN_684; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_686 = 4'hd == _T_401 ? csrExceptionVec_13 : _GEN_685; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_687 = 4'he == _T_401 ? 1'h0 : _GEN_686; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_688 = 4'hf == _T_401 ? csrExceptionVec_15 : _GEN_687; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_402 = _GEN_688 ? _T_401 : 4'h2; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_691 = 4'h2 == _T_402 ? csrExceptionVec_2 : 4'h1 == _T_402 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_692 = 4'h3 == _T_402 ? csrExceptionVec_3 : _GEN_691; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_693 = 4'h4 == _T_402 ? io_cfIn_exceptionVec_4 : _GEN_692; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_694 = 4'h5 == _T_402 ? 1'h0 : _GEN_693; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_695 = 4'h6 == _T_402 ? io_cfIn_exceptionVec_6 : _GEN_694; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_696 = 4'h7 == _T_402 ? 1'h0 : _GEN_695; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_697 = 4'h8 == _T_402 ? csrExceptionVec_8 : _GEN_696; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_698 = 4'h9 == _T_402 ? csrExceptionVec_9 : _GEN_697; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_699 = 4'ha == _T_402 ? 1'h0 : _GEN_698; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_700 = 4'hb == _T_402 ? csrExceptionVec_11 : _GEN_699; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_701 = 4'hc == _T_402 ? io_cfIn_exceptionVec_12 : _GEN_700; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_702 = 4'hd == _T_402 ? csrExceptionVec_13 : _GEN_701; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_703 = 4'he == _T_402 ? 1'h0 : _GEN_702; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_704 = 4'hf == _T_402 ? csrExceptionVec_15 : _GEN_703; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_403 = _GEN_704 ? _T_402 : 4'h0; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_707 = 4'h2 == _T_403 ? csrExceptionVec_2 : 4'h1 == _T_403 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_708 = 4'h3 == _T_403 ? csrExceptionVec_3 : _GEN_707; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_709 = 4'h4 == _T_403 ? io_cfIn_exceptionVec_4 : _GEN_708; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_710 = 4'h5 == _T_403 ? 1'h0 : _GEN_709; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_711 = 4'h6 == _T_403 ? io_cfIn_exceptionVec_6 : _GEN_710; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_712 = 4'h7 == _T_403 ? 1'h0 : _GEN_711; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_713 = 4'h8 == _T_403 ? csrExceptionVec_8 : _GEN_712; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_714 = 4'h9 == _T_403 ? csrExceptionVec_9 : _GEN_713; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_715 = 4'ha == _T_403 ? 1'h0 : _GEN_714; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_716 = 4'hb == _T_403 ? csrExceptionVec_11 : _GEN_715; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_717 = 4'hc == _T_403 ? io_cfIn_exceptionVec_12 : _GEN_716; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_718 = 4'hd == _T_403 ? csrExceptionVec_13 : _GEN_717; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_719 = 4'he == _T_403 ? 1'h0 : _GEN_718; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_720 = 4'hf == _T_403 ? csrExceptionVec_15 : _GEN_719; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_404 = _GEN_720 ? _T_403 : 4'hb; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_723 = 4'h2 == _T_404 ? csrExceptionVec_2 : 4'h1 == _T_404 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_724 = 4'h3 == _T_404 ? csrExceptionVec_3 : _GEN_723; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_725 = 4'h4 == _T_404 ? io_cfIn_exceptionVec_4 : _GEN_724; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_726 = 4'h5 == _T_404 ? 1'h0 : _GEN_725; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_727 = 4'h6 == _T_404 ? io_cfIn_exceptionVec_6 : _GEN_726; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_728 = 4'h7 == _T_404 ? 1'h0 : _GEN_727; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_729 = 4'h8 == _T_404 ? csrExceptionVec_8 : _GEN_728; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_730 = 4'h9 == _T_404 ? csrExceptionVec_9 : _GEN_729; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_731 = 4'ha == _T_404 ? 1'h0 : _GEN_730; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_732 = 4'hb == _T_404 ? csrExceptionVec_11 : _GEN_731; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_733 = 4'hc == _T_404 ? io_cfIn_exceptionVec_12 : _GEN_732; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_734 = 4'hd == _T_404 ? csrExceptionVec_13 : _GEN_733; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_735 = 4'he == _T_404 ? 1'h0 : _GEN_734; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_736 = 4'hf == _T_404 ? csrExceptionVec_15 : _GEN_735; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_405 = _GEN_736 ? _T_404 : 4'h9; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_739 = 4'h2 == _T_405 ? csrExceptionVec_2 : 4'h1 == _T_405 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_740 = 4'h3 == _T_405 ? csrExceptionVec_3 : _GEN_739; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_741 = 4'h4 == _T_405 ? io_cfIn_exceptionVec_4 : _GEN_740; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_742 = 4'h5 == _T_405 ? 1'h0 : _GEN_741; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_743 = 4'h6 == _T_405 ? io_cfIn_exceptionVec_6 : _GEN_742; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_744 = 4'h7 == _T_405 ? 1'h0 : _GEN_743; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_745 = 4'h8 == _T_405 ? csrExceptionVec_8 : _GEN_744; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_746 = 4'h9 == _T_405 ? csrExceptionVec_9 : _GEN_745; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_747 = 4'ha == _T_405 ? 1'h0 : _GEN_746; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_748 = 4'hb == _T_405 ? csrExceptionVec_11 : _GEN_747; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_749 = 4'hc == _T_405 ? io_cfIn_exceptionVec_12 : _GEN_748; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_750 = 4'hd == _T_405 ? csrExceptionVec_13 : _GEN_749; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_751 = 4'he == _T_405 ? 1'h0 : _GEN_750; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_752 = 4'hf == _T_405 ? csrExceptionVec_15 : _GEN_751; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_406 = _GEN_752 ? _T_405 : 4'h8; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_755 = 4'h2 == _T_406 ? csrExceptionVec_2 : 4'h1 == _T_406 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_756 = 4'h3 == _T_406 ? csrExceptionVec_3 : _GEN_755; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_757 = 4'h4 == _T_406 ? io_cfIn_exceptionVec_4 : _GEN_756; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_758 = 4'h5 == _T_406 ? 1'h0 : _GEN_757; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_759 = 4'h6 == _T_406 ? io_cfIn_exceptionVec_6 : _GEN_758; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_760 = 4'h7 == _T_406 ? 1'h0 : _GEN_759; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_761 = 4'h8 == _T_406 ? csrExceptionVec_8 : _GEN_760; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_762 = 4'h9 == _T_406 ? csrExceptionVec_9 : _GEN_761; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_763 = 4'ha == _T_406 ? 1'h0 : _GEN_762; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_764 = 4'hb == _T_406 ? csrExceptionVec_11 : _GEN_763; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_765 = 4'hc == _T_406 ? io_cfIn_exceptionVec_12 : _GEN_764; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_766 = 4'hd == _T_406 ? csrExceptionVec_13 : _GEN_765; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_767 = 4'he == _T_406 ? 1'h0 : _GEN_766; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_768 = 4'hf == _T_406 ? csrExceptionVec_15 : _GEN_767; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_407 = _GEN_768 ? _T_406 : 4'h6; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_771 = 4'h2 == _T_407 ? csrExceptionVec_2 : 4'h1 == _T_407 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_772 = 4'h3 == _T_407 ? csrExceptionVec_3 : _GEN_771; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_773 = 4'h4 == _T_407 ? io_cfIn_exceptionVec_4 : _GEN_772; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_774 = 4'h5 == _T_407 ? 1'h0 : _GEN_773; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_775 = 4'h6 == _T_407 ? io_cfIn_exceptionVec_6 : _GEN_774; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_776 = 4'h7 == _T_407 ? 1'h0 : _GEN_775; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_777 = 4'h8 == _T_407 ? csrExceptionVec_8 : _GEN_776; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_778 = 4'h9 == _T_407 ? csrExceptionVec_9 : _GEN_777; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_779 = 4'ha == _T_407 ? 1'h0 : _GEN_778; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_780 = 4'hb == _T_407 ? csrExceptionVec_11 : _GEN_779; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_781 = 4'hc == _T_407 ? io_cfIn_exceptionVec_12 : _GEN_780; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_782 = 4'hd == _T_407 ? csrExceptionVec_13 : _GEN_781; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_783 = 4'he == _T_407 ? 1'h0 : _GEN_782; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_784 = 4'hf == _T_407 ? csrExceptionVec_15 : _GEN_783; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_408 = _GEN_784 ? _T_407 : 4'h4; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_787 = 4'h2 == _T_408 ? csrExceptionVec_2 : 4'h1 == _T_408 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_788 = 4'h3 == _T_408 ? csrExceptionVec_3 : _GEN_787; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_789 = 4'h4 == _T_408 ? io_cfIn_exceptionVec_4 : _GEN_788; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_790 = 4'h5 == _T_408 ? 1'h0 : _GEN_789; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_791 = 4'h6 == _T_408 ? io_cfIn_exceptionVec_6 : _GEN_790; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_792 = 4'h7 == _T_408 ? 1'h0 : _GEN_791; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_793 = 4'h8 == _T_408 ? csrExceptionVec_8 : _GEN_792; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_794 = 4'h9 == _T_408 ? csrExceptionVec_9 : _GEN_793; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_795 = 4'ha == _T_408 ? 1'h0 : _GEN_794; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_796 = 4'hb == _T_408 ? csrExceptionVec_11 : _GEN_795; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_797 = 4'hc == _T_408 ? io_cfIn_exceptionVec_12 : _GEN_796; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_798 = 4'hd == _T_408 ? csrExceptionVec_13 : _GEN_797; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_799 = 4'he == _T_408 ? 1'h0 : _GEN_798; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_800 = 4'hf == _T_408 ? csrExceptionVec_15 : _GEN_799; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_409 = _GEN_800 ? _T_408 : 4'hf; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_803 = 4'h2 == _T_409 ? csrExceptionVec_2 : 4'h1 == _T_409 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_804 = 4'h3 == _T_409 ? csrExceptionVec_3 : _GEN_803; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_805 = 4'h4 == _T_409 ? io_cfIn_exceptionVec_4 : _GEN_804; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_806 = 4'h5 == _T_409 ? 1'h0 : _GEN_805; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_807 = 4'h6 == _T_409 ? io_cfIn_exceptionVec_6 : _GEN_806; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_808 = 4'h7 == _T_409 ? 1'h0 : _GEN_807; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_809 = 4'h8 == _T_409 ? csrExceptionVec_8 : _GEN_808; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_810 = 4'h9 == _T_409 ? csrExceptionVec_9 : _GEN_809; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_811 = 4'ha == _T_409 ? 1'h0 : _GEN_810; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_812 = 4'hb == _T_409 ? csrExceptionVec_11 : _GEN_811; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_813 = 4'hc == _T_409 ? io_cfIn_exceptionVec_12 : _GEN_812; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_814 = 4'hd == _T_409 ? csrExceptionVec_13 : _GEN_813; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_815 = 4'he == _T_409 ? 1'h0 : _GEN_814; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_816 = 4'hf == _T_409 ? csrExceptionVec_15 : _GEN_815; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_410 = _GEN_816 ? _T_409 : 4'hd; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_819 = 4'h2 == _T_410 ? csrExceptionVec_2 : 4'h1 == _T_410 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_820 = 4'h3 == _T_410 ? csrExceptionVec_3 : _GEN_819; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_821 = 4'h4 == _T_410 ? io_cfIn_exceptionVec_4 : _GEN_820; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_822 = 4'h5 == _T_410 ? 1'h0 : _GEN_821; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_823 = 4'h6 == _T_410 ? io_cfIn_exceptionVec_6 : _GEN_822; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_824 = 4'h7 == _T_410 ? 1'h0 : _GEN_823; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_825 = 4'h8 == _T_410 ? csrExceptionVec_8 : _GEN_824; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_826 = 4'h9 == _T_410 ? csrExceptionVec_9 : _GEN_825; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_827 = 4'ha == _T_410 ? 1'h0 : _GEN_826; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_828 = 4'hb == _T_410 ? csrExceptionVec_11 : _GEN_827; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_829 = 4'hc == _T_410 ? io_cfIn_exceptionVec_12 : _GEN_828; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_830 = 4'hd == _T_410 ? csrExceptionVec_13 : _GEN_829; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_831 = 4'he == _T_410 ? 1'h0 : _GEN_830; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_832 = 4'hf == _T_410 ? csrExceptionVec_15 : _GEN_831; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] _T_411 = _GEN_832 ? _T_410 : 4'h7; // @[SIMD_CSR.scala 809:68]
  wire  _GEN_835 = 4'h2 == _T_411 ? csrExceptionVec_2 : 4'h1 == _T_411 & io_cfIn_exceptionVec_1; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_836 = 4'h3 == _T_411 ? csrExceptionVec_3 : _GEN_835; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_837 = 4'h4 == _T_411 ? io_cfIn_exceptionVec_4 : _GEN_836; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_838 = 4'h5 == _T_411 ? 1'h0 : _GEN_837; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_839 = 4'h6 == _T_411 ? io_cfIn_exceptionVec_6 : _GEN_838; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_840 = 4'h7 == _T_411 ? 1'h0 : _GEN_839; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_841 = 4'h8 == _T_411 ? csrExceptionVec_8 : _GEN_840; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_842 = 4'h9 == _T_411 ? csrExceptionVec_9 : _GEN_841; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_843 = 4'ha == _T_411 ? 1'h0 : _GEN_842; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_844 = 4'hb == _T_411 ? csrExceptionVec_11 : _GEN_843; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_845 = 4'hc == _T_411 ? io_cfIn_exceptionVec_12 : _GEN_844; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_846 = 4'hd == _T_411 ? csrExceptionVec_13 : _GEN_845; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_847 = 4'he == _T_411 ? 1'h0 : _GEN_846; // @[SIMD_CSR.scala 809:{68,68}]
  wire  _GEN_848 = 4'hf == _T_411 ? csrExceptionVec_15 : _GEN_847; // @[SIMD_CSR.scala 809:{68,68}]
  wire [3:0] exceptionNO = _GEN_848 ? _T_411 : 4'h5; // @[SIMD_CSR.scala 809:68]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid & _T_55; // @[SIMD_CSR.scala 812:75]
  wire [63:0] _T_416 = {raiseIntr,63'h0}; // @[Cat.scala 30:58]
  wire [3:0] _T_417 = raiseIntr ? intrNO : exceptionNO; // @[SIMD_CSR.scala 813:54]
  wire [63:0] _GEN_934 = {{60'd0}, _T_417}; // @[SIMD_CSR.scala 813:49]
  wire [63:0] causeNO = _T_416 | _GEN_934; // @[SIMD_CSR.scala 813:49]
  wire [63:0] _T_483 = raiseIntr ? mideleg : medeleg; // @[SIMD_CSR.scala 823:20]
  wire [63:0] _T_485 = _T_483 >> causeNO[3:0]; // @[SIMD_CSR.scala 823:50]
  wire  delegS = _T_485[0] & _T_247; // @[SIMD_CSR.scala 823:66]
  wire  _T_489 = io_cfIn_exceptionVec_12 | csrExceptionVec_13 | csrExceptionVec_15; // @[SIMD_CSR.scala 826:88]
  wire  _T_490 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[SIMD_CSR.scala 827:58]
  wire [24:0] _T_493 = LSUADDR[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_494 = {_T_493,LSUADDR[38:0]}; // @[Cat.scala 30:58]
  wire [38:0] _T_496 = io_cfIn_pc + 39'h2; // @[SIMD_CSR.scala 836:109]
  wire [24:0] _T_500 = _T_496[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_501 = {_T_500,_T_496}; // @[Cat.scala 30:58]
  wire [24:0] _T_505 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_506 = {_T_505,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_507 = io_cfIn_crossPageIPFFix ? _T_501 : _T_506; // @[SIMD_CSR.scala 836:63]
  wire [24:0] _T_510 = io_dmemMMU_addr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_511 = {_T_510,io_dmemMMU_addr}; // @[Cat.scala 30:58]
  wire [63:0] _T_512 = io_cfIn_exceptionVec_12 ? _T_507 : _T_511; // @[SIMD_CSR.scala 836:26]
  wire [63:0] _T_513 = _T_490 ? _T_494 : _T_512; // @[SIMD_CSR.scala 835:23]
  wire [1:0] _GEN_853 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[SIMD_CSR.scala 837:19 840:22]
  wire  _GEN_854 = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[SIMD_CSR.scala 837:19 841:24]
  wire  _GEN_855 = delegS ? 1'h0 : mstatusStruct_ie_s; // @[SIMD_CSR.scala 837:19 842:23]
  wire [38:0] _GEN_858 = delegS ? stvec[38:0] : mtvec[38:0]; // @[SIMD_CSR.scala 837:19 849:18 862:18]
  wire [1:0] _GEN_861 = delegS ? mstatusStruct_mpp : priviledgeMode; // @[SIMD_CSR.scala 837:19 853:22]
  wire  _GEN_862 = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[SIMD_CSR.scala 837:19 854:24]
  wire  _GEN_863 = delegS & mstatusStruct_ie_m; // @[SIMD_CSR.scala 837:19 855:23]
  wire  _GEN_870 = isSret ? mstatusStruct_pie_s : mstatusStruct_ie_s; // @[SIMD_CSR.scala 873:25 875:23]
  wire  _GEN_881 = isMret ? mstatusStruct_ie_s : _GEN_870; // @[SIMD_CSR.scala 867:19]
  wire  _GEN_891 = isRet ? _GEN_881 : mstatusStruct_ie_s; // @[SIMD_CSR.scala 866:20]
  wire  mstatusNew_ie_s = raiseExceptionIntr ? _GEN_855 : _GEN_891; // @[SIMD_CSR.scala 825:29]
  wire  _GEN_866 = isUret ? mstatusStruct_pie_u : mstatusStruct_ie_u; // @[SIMD_CSR.scala 879:25 881:23]
  wire  _GEN_874 = isSret ? mstatusStruct_ie_u : _GEN_866; // @[SIMD_CSR.scala 873:25]
  wire  _GEN_884 = isMret ? mstatusStruct_ie_u : _GEN_874; // @[SIMD_CSR.scala 867:19]
  wire  _GEN_894 = isRet ? _GEN_884 : mstatusStruct_ie_u; // @[SIMD_CSR.scala 866:20]
  wire  mstatusNew_ie_u = raiseExceptionIntr ? mstatusStruct_ie_u : _GEN_894; // @[SIMD_CSR.scala 825:29]
  wire  _GEN_871 = isSret | mstatusStruct_pie_s; // @[SIMD_CSR.scala 873:25 876:24]
  wire  _GEN_882 = isMret ? mstatusStruct_pie_s : _GEN_871; // @[SIMD_CSR.scala 867:19]
  wire  _GEN_892 = isRet ? _GEN_882 : mstatusStruct_pie_s; // @[SIMD_CSR.scala 866:20]
  wire  mstatusNew_pie_s = raiseExceptionIntr ? _GEN_854 : _GEN_892; // @[SIMD_CSR.scala 825:29]
  wire  _GEN_867 = isUret | mstatusStruct_pie_u; // @[SIMD_CSR.scala 879:25 882:24]
  wire  _GEN_875 = isSret ? mstatusStruct_pie_u : _GEN_867; // @[SIMD_CSR.scala 873:25]
  wire  _GEN_885 = isMret ? mstatusStruct_pie_u : _GEN_875; // @[SIMD_CSR.scala 867:19]
  wire  _GEN_895 = isRet ? _GEN_885 : mstatusStruct_pie_u; // @[SIMD_CSR.scala 866:20]
  wire  mstatusNew_pie_u = raiseExceptionIntr ? mstatusStruct_pie_u : _GEN_895; // @[SIMD_CSR.scala 825:29]
  wire  _GEN_877 = isMret ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[SIMD_CSR.scala 867:19 869:23]
  wire  _GEN_887 = isRet ? _GEN_877 : mstatusStruct_ie_m; // @[SIMD_CSR.scala 866:20]
  wire  mstatusNew_ie_m = raiseExceptionIntr ? _GEN_863 : _GEN_887; // @[SIMD_CSR.scala 825:29]
  wire [5:0] lo_lo_12 = {mstatusNew_pie_s,mstatusNew_pie_u,mstatusNew_ie_m,mstatusStruct_ie_h,mstatusNew_ie_s,
    mstatusNew_ie_u}; // @[SIMD_CSR.scala 864:27]
  wire  _GEN_872 = isSret ? 1'h0 : mstatusStruct_spp; // @[SIMD_CSR.scala 873:25 877:22]
  wire  _GEN_883 = isMret ? mstatusStruct_spp : _GEN_872; // @[SIMD_CSR.scala 867:19]
  wire  _GEN_893 = isRet ? _GEN_883 : mstatusStruct_spp; // @[SIMD_CSR.scala 866:20]
  wire [1:0] _GEN_900 = raiseExceptionIntr ? _GEN_853 : {{1'd0}, _GEN_893}; // @[SIMD_CSR.scala 825:29]
  wire  mstatusNew_spp = _GEN_900[0];
  wire  _GEN_878 = isMret | mstatusStruct_pie_m; // @[SIMD_CSR.scala 867:19 870:24]
  wire  _GEN_888 = isRet ? _GEN_878 : mstatusStruct_pie_m; // @[SIMD_CSR.scala 866:20]
  wire  mstatusNew_pie_m = raiseExceptionIntr ? _GEN_862 : _GEN_888; // @[SIMD_CSR.scala 825:29]
  wire [1:0] _GEN_879 = isMret ? 2'h0 : mstatusStruct_mpp; // @[SIMD_CSR.scala 867:19 871:22]
  wire [1:0] _GEN_889 = isRet ? _GEN_879 : mstatusStruct_mpp; // @[SIMD_CSR.scala 866:20]
  wire [1:0] mstatusNew_mpp = raiseExceptionIntr ? _GEN_861 : _GEN_889; // @[SIMD_CSR.scala 825:29]
  wire [14:0] lo_12 = {mstatusStruct_fs,mstatusNew_mpp,mstatusStruct_hpp,mstatusNew_spp,mstatusNew_pie_m,
    mstatusStruct_pie_h,lo_lo_12}; // @[SIMD_CSR.scala 864:27]
  wire [6:0] hi_lo_12 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,
    mstatusStruct_xs}; // @[SIMD_CSR.scala 864:27]
  wire [63:0] _T_574 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_12,lo_12}; // @[SIMD_CSR.scala 864:27]
  wire [1:0] _T_576 = {1'h0,mstatusStruct_spp}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_865 = isUret ? 2'h0 : priviledgeMode; // @[SIMD_CSR.scala 879:25 880:22 638:31]
  wire [1:0] _GEN_869 = isSret ? _T_576 : _GEN_865; // @[SIMD_CSR.scala 873:25 874:22]
  wire [38:0] _GEN_873 = isSret ? sepc[38:0] : 39'h0; // @[SIMD_CSR.scala 873:25 878:17]
  wire [38:0] _GEN_880 = isMret ? mepc[38:0] : _GEN_873; // @[SIMD_CSR.scala 867:19 872:17]
  wire [38:0] _GEN_890 = isRet ? _GEN_880 : 39'h0; // @[SIMD_CSR.scala 866:20]
  wire [38:0] trapTarget = raiseExceptionIntr ? _GEN_858 : 39'h0; // @[SIMD_CSR.scala 825:29]
  wire [38:0] retTarget = raiseExceptionIntr ? 39'h0 : _GEN_890; // @[SIMD_CSR.scala 825:29]
  wire [38:0] _T_594 = io_cfIn_pc + 39'h4; // @[SIMD_CSR.scala 918:60]
  wire [38:0] _T_595 = raiseExceptionIntr ? trapTarget : retTarget; // @[SIMD_CSR.scala 918:70]
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1 & io_ctrlIn_isMou; // @[SIMD_CSR.scala 921:58]
  wire  flushTLB = io_in_valid & _T_58 & io_ctrlIn_isMou; // @[SIMD_CSR.scala 925:59]
  assign io_out_bits = addr == 12'h100 ? _T_70 : _GEN_512; // @[SIMD_CSR.scala 662:27 663:11]
  assign io_redirect_target = resetSatp | io_ctrlIn_isMou ? _T_594 : _T_595; // @[SIMD_CSR.scala 918:28]
  assign io_redirect_valid = io_in_valid & (JumpType | io_ctrlIn_isMou) | raiseExceptionIntr | resetSatp; // @[SIMD_CSR.scala 916:77]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[SIMD_CSR.scala 904:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[SIMD_CSR.scala 905:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[SIMD_CSR.scala 599:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[SIMD_CSR.scala 599:39]
  assign io_wenFix = raiseException & io_in_valid & _T_55; // @[SIMD_CSR.scala 915:40]
  assign flushICache_0 = flushICache;
  assign satp_0 = satp;
  assign lr_0 = lr;
  assign intrVec_0 = intrVec;
  assign flushTLB_0 = flushTLB;
  assign lrAddr_0 = lrAddr;
  always @(posedge clock) begin
    if (reset) begin // @[SIMD_CSR.scala 560:19]
      lr <= 1'h0; // @[SIMD_CSR.scala 560:19]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      lr <= 1'h0; // @[SIMD_CSR.scala 865:8]
    end else if (isRet) begin // @[SIMD_CSR.scala 866:20]
      lr <= 1'h0; // @[SIMD_CSR.scala 886:7]
    end else if (set_lr) begin // @[SIMD_CSR.scala 568:14]
      lr <= set_lr_val; // @[SIMD_CSR.scala 569:8]
    end
    if (reset) begin // @[SIMD_CSR.scala 561:23]
      lrAddr <= 64'h0; // @[SIMD_CSR.scala 561:23]
    end else if (set_lr) begin // @[SIMD_CSR.scala 568:14]
      lrAddr <= set_lr_addr; // @[SIMD_CSR.scala 570:12]
    end
    if (reset) begin // @[SIMD_CSR.scala 575:22]
      mtvec <= 64'h0; // @[SIMD_CSR.scala 575:22]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          mtvec <= _GEN_465;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 576:27]
      mcounteren <= 64'h0; // @[SIMD_CSR.scala 576:27]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          mcounteren <= _GEN_466;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 577:23]
      mcause <= 64'h0; // @[SIMD_CSR.scala 577:23]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        mcause <= _GEN_559;
      end else begin
        mcause <= causeNO; // @[SIMD_CSR.scala 851:14]
      end
    end else begin
      mcause <= _GEN_559;
    end
    if (reset) begin // @[SIMD_CSR.scala 578:22]
      mtval <= 64'h0; // @[SIMD_CSR.scala 578:22]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        mtval <= _GEN_560;
      end else if (_T_489 | _T_490) begin // @[SIMD_CSR.scala 844:38]
        mtval <= _T_513; // @[SIMD_CSR.scala 845:15]
      end else begin
        mtval <= 64'h0; // @[SIMD_CSR.scala 847:15]
      end
    end else begin
      mtval <= _GEN_560;
    end
    if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        mepc <= _GEN_558;
      end else begin
        mepc <= _T_506; // @[SIMD_CSR.scala 852:12]
      end
    end else begin
      mepc <= _GEN_558;
    end
    if (reset) begin // @[SIMD_CSR.scala 581:20]
      mie <= 64'h0; // @[SIMD_CSR.scala 581:20]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (addr == 12'h104) begin // @[SIMD_CSR.scala 666:29]
        if (RegWen & io_cfIn_pc != 39'h80001f04) begin // @[SIMD_CSR.scala 668:49]
          mie <= _T_109; // @[SIMD_CSR.scala 668:54]
        end
      end else if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
        mie <= _GEN_464;
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 583:24]
      mipReg <= 64'h0; // @[SIMD_CSR.scala 583:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          mipReg <= _GEN_480;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 598:24]
      mstatus <= 64'h1800; // @[SIMD_CSR.scala 598:24]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      mstatus <= _T_574; // @[SIMD_CSR.scala 864:13]
    end else if (isRet) begin // @[SIMD_CSR.scala 866:20]
      mstatus <= _T_574; // @[SIMD_CSR.scala 885:13]
    end else if (addr == 12'h100) begin // @[SIMD_CSR.scala 662:27]
      mstatus <= _GEN_2;
    end else begin
      mstatus <= _GEN_522;
    end
    if (reset) begin // @[SIMD_CSR.scala 600:24]
      medeleg <= 64'h0; // @[SIMD_CSR.scala 600:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          medeleg <= _GEN_462;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 601:24]
      mideleg <= 64'h0; // @[SIMD_CSR.scala 601:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          mideleg <= _GEN_463;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 602:25]
      mscratch <= 64'h0; // @[SIMD_CSR.scala 602:25]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          mscratch <= _GEN_467;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 604:24]
      pmpcfg0 <= 64'h0; // @[SIMD_CSR.scala 604:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpcfg0 <= _GEN_471;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 605:24]
      pmpcfg1 <= 64'h0; // @[SIMD_CSR.scala 605:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpcfg1 <= _GEN_472;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 606:24]
      pmpcfg2 <= 64'h0; // @[SIMD_CSR.scala 606:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpcfg2 <= _GEN_473;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 607:24]
      pmpcfg3 <= 64'h0; // @[SIMD_CSR.scala 607:24]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpcfg3 <= _GEN_474;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 608:25]
      pmpaddr0 <= 64'h0; // @[SIMD_CSR.scala 608:25]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpaddr0 <= _GEN_475;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 609:25]
      pmpaddr1 <= 64'h0; // @[SIMD_CSR.scala 609:25]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpaddr1 <= _GEN_476;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 610:25]
      pmpaddr2 <= 64'h0; // @[SIMD_CSR.scala 610:25]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpaddr2 <= _GEN_477;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 611:25]
      pmpaddr3 <= 64'h0; // @[SIMD_CSR.scala 611:25]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          pmpaddr3 <= _GEN_478;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 613:22]
      vxsat <= 64'h0; // @[SIMD_CSR.scala 613:22]
    end else if (OVWEN_0) begin // @[SIMD_CSR.scala 775:14]
      vxsat <= 64'h1; // @[SIMD_CSR.scala 775:21]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        vxsat <= _GEN_509;
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 620:22]
      stvec <= 64'h0; // @[SIMD_CSR.scala 620:22]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (addr == 12'h105) begin // @[SIMD_CSR.scala 669:31]
          stvec <= _GEN_4;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 623:21]
      satp <= 64'h0; // @[SIMD_CSR.scala 623:21]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          satp <= _GEN_459;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 624:21]
      sepc <= 64'h0; // @[SIMD_CSR.scala 624:21]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        sepc <= _T_506; // @[SIMD_CSR.scala 839:12]
      end else begin
        sepc <= _GEN_548;
      end
    end else begin
      sepc <= _GEN_548;
    end
    if (reset) begin // @[SIMD_CSR.scala 625:23]
      scause <= 64'h0; // @[SIMD_CSR.scala 625:23]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        scause <= causeNO; // @[SIMD_CSR.scala 838:14]
      end else begin
        scause <= _GEN_549;
      end
    end else begin
      scause <= _GEN_549;
    end
    if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        if (_T_489 | _T_490) begin // @[SIMD_CSR.scala 844:38]
          if (_T_490) begin // @[SIMD_CSR.scala 835:23]
            stval <= _T_494;
          end else begin
            stval <= _T_512;
          end
        end else begin
          stval <= 64'h0; // @[SIMD_CSR.scala 847:15]
        end
      end else begin
        stval <= _GEN_550;
      end
    end else begin
      stval <= _GEN_550;
    end
    if (reset) begin // @[SIMD_CSR.scala 627:25]
      sscratch <= 64'h0; // @[SIMD_CSR.scala 627:25]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          sscratch <= _GEN_455;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 628:27]
      scounteren <= 64'h0; // @[SIMD_CSR.scala 628:27]
    end else if (!(addr == 12'h100)) begin // @[SIMD_CSR.scala 662:27]
      if (!(addr == 12'h104)) begin // @[SIMD_CSR.scala 666:29]
        if (!(addr == 12'h105)) begin // @[SIMD_CSR.scala 669:31]
          scounteren <= _GEN_454;
        end
      end
    end
    if (reset) begin // @[SIMD_CSR.scala 638:31]
      priviledgeMode <= 2'h3; // @[SIMD_CSR.scala 638:31]
    end else if (raiseExceptionIntr) begin // @[SIMD_CSR.scala 825:29]
      if (delegS) begin // @[SIMD_CSR.scala 837:19]
        priviledgeMode <= 2'h1; // @[SIMD_CSR.scala 843:22]
      end else begin
        priviledgeMode <= 2'h3; // @[SIMD_CSR.scala 856:22]
      end
    end else if (isRet) begin // @[SIMD_CSR.scala 866:20]
      if (isMret) begin // @[SIMD_CSR.scala 867:19]
        priviledgeMode <= mstatusStruct_mpp; // @[SIMD_CSR.scala 868:22]
      end else begin
        priviledgeMode <= _GEN_869;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lr = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  lrAddr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mtvec = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcounteren = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mcause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mtval = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mepc = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mie = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mipReg = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  mstatus = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  medeleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mideleg = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  mscratch = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg0 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg1 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg2 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpcfg3 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr0 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr1 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr2 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  pmpaddr3 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  vxsat = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  stvec = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  satp = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  sepc = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  scause = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  stval = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  sscratch = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  scounteren = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  priviledgeMode = _RAND_29[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PerfU(
  input         clock,
  input         reset,
  input         perfCntCondMultiCommit3,
  input         perfCntCondMultiCommit6,
  output [63:0] perfCnts_2_0,
  input         perfCntCondMinstret,
  input         perfCntCondMultiCommit2,
  input         perfCntCondMultiCommit5,
  input         perfCntCondMultiCommit4,
  input         perfCntCondMultiCommit
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] perfCnts_2; // @[PerfU.scala 14:47]
  wire  _WIRE = 1'h1;
  wire [63:0] _T_11 = perfCnts_2 + 64'h1; // @[PerfU.scala 64:71]
  wire [63:0] _GEN_2 = perfCntCondMinstret ? _T_11 : perfCnts_2; // @[PerfU.scala 14:47 64:{62,66}]
  wire [63:0] _T_13 = perfCnts_2 + 64'h2; // @[PerfU.scala 73:88]
  wire [63:0] _T_15 = perfCnts_2 + 64'h3; // @[PerfU.scala 75:88]
  wire [63:0] _T_17 = perfCnts_2 + 64'h4; // @[PerfU.scala 77:88]
  wire [63:0] _T_19 = perfCnts_2 + 64'h5; // @[PerfU.scala 79:88]
  wire [63:0] _T_21 = perfCnts_2 + 64'h6; // @[PerfU.scala 81:88]
  wire [63:0] _GEN_3 = perfCntCondMultiCommit6 ? _T_21 : _GEN_2; // @[PerfU.scala 80:72 81:62]
  wire [63:0] _GEN_4 = perfCntCondMultiCommit5 ? _T_19 : _GEN_3; // @[PerfU.scala 78:72 79:62]
  wire [63:0] _GEN_5 = perfCntCondMultiCommit4 ? _T_17 : _GEN_4; // @[PerfU.scala 76:72 77:62]
  assign perfCnts_2_0 = perfCnts_2;
  always @(posedge clock) begin
    if (reset) begin // @[PerfU.scala 14:47]
      perfCnts_2 <= 64'h0; // @[PerfU.scala 14:47]
    end else if (perfCntCondMultiCommit) begin // @[PerfU.scala 72:35]
      if (perfCntCondMultiCommit2) begin // @[PerfU.scala 72:68]
        perfCnts_2 <= _T_13; // @[PerfU.scala 73:62]
      end else if (perfCntCondMultiCommit3) begin // @[PerfU.scala 74:72]
        perfCnts_2 <= _T_15; // @[PerfU.scala 75:62]
      end else begin
        perfCnts_2 <= _GEN_5;
      end
    end else if (perfCntCondMinstret) begin // @[PerfU.scala 64:62]
      perfCnts_2 <= _T_11; // @[PerfU.scala 64:66]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  perfCnts_2 = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module new_SIMD_EXU(
  input         clock,
  input         reset,
  output        io__in_0_ready,
  input         io__in_0_valid,
  input  [63:0] io__in_0_bits_cf_instr,
  input  [38:0] io__in_0_bits_cf_pc,
  input  [38:0] io__in_0_bits_cf_pnpc,
  input  [3:0]  io__in_0_bits_cf_brIdx,
  input  [63:0] io__in_0_bits_cf_runahead_checkpoint_id,
  input  [6:0]  io__in_0_bits_ctrl_fuOpType,
  input         io__in_0_bits_ctrl_rfWen,
  input  [4:0]  io__in_0_bits_ctrl_rfDest,
  input  [63:0] io__in_0_bits_data_src1,
  input  [63:0] io__in_0_bits_data_src2,
  input  [63:0] io__in_0_bits_data_imm,
  input  [4:0]  io__in_0_bits_InstNo,
  input         io__in_0_bits_InstFlag,
  output        io__in_1_ready,
  input         io__in_1_valid,
  input  [38:0] io__in_1_bits_cf_pc,
  input         io__in_1_bits_cf_exceptionVec_1,
  input         io__in_1_bits_cf_exceptionVec_2,
  input         io__in_1_bits_cf_exceptionVec_12,
  input         io__in_1_bits_cf_intrVec_0,
  input         io__in_1_bits_cf_intrVec_1,
  input         io__in_1_bits_cf_intrVec_2,
  input         io__in_1_bits_cf_intrVec_3,
  input         io__in_1_bits_cf_intrVec_4,
  input         io__in_1_bits_cf_intrVec_5,
  input         io__in_1_bits_cf_intrVec_6,
  input         io__in_1_bits_cf_intrVec_7,
  input         io__in_1_bits_cf_intrVec_8,
  input         io__in_1_bits_cf_intrVec_9,
  input         io__in_1_bits_cf_intrVec_10,
  input         io__in_1_bits_cf_intrVec_11,
  input         io__in_1_bits_cf_crossPageIPFFix,
  input  [63:0] io__in_1_bits_cf_runahead_checkpoint_id,
  input  [6:0]  io__in_1_bits_ctrl_fuOpType,
  input         io__in_1_bits_ctrl_rfWen,
  input  [4:0]  io__in_1_bits_ctrl_rfDest,
  input         io__in_1_bits_ctrl_isMou,
  input  [63:0] io__in_1_bits_data_src1,
  input  [63:0] io__in_1_bits_data_src2,
  input  [4:0]  io__in_1_bits_InstNo,
  input         io__in_1_bits_InstFlag,
  output        io__in_2_ready,
  input         io__in_2_valid,
  input  [63:0] io__in_2_bits_cf_instr,
  input  [38:0] io__in_2_bits_cf_pc,
  input  [63:0] io__in_2_bits_cf_runahead_checkpoint_id,
  input  [4:0]  io__in_2_bits_cf_instrType,
  input  [6:0]  io__in_2_bits_ctrl_fuOpType,
  input  [2:0]  io__in_2_bits_ctrl_funct3,
  input         io__in_2_bits_ctrl_func24,
  input         io__in_2_bits_ctrl_func23,
  input         io__in_2_bits_ctrl_rfWen,
  input  [4:0]  io__in_2_bits_ctrl_rfDest,
  input  [63:0] io__in_2_bits_data_src1,
  input  [63:0] io__in_2_bits_data_src2,
  input  [63:0] io__in_2_bits_data_src3,
  input  [4:0]  io__in_2_bits_InstNo,
  input         io__in_2_bits_InstFlag,
  output        io__in_3_ready,
  input         io__in_3_valid,
  input  [63:0] io__in_3_bits_cf_instr,
  input  [38:0] io__in_3_bits_cf_pc,
  input  [63:0] io__in_3_bits_cf_runahead_checkpoint_id,
  input  [4:0]  io__in_3_bits_cf_instrType,
  input  [6:0]  io__in_3_bits_ctrl_fuOpType,
  input  [2:0]  io__in_3_bits_ctrl_funct3,
  input         io__in_3_bits_ctrl_func24,
  input         io__in_3_bits_ctrl_func23,
  input         io__in_3_bits_ctrl_rfWen,
  input  [4:0]  io__in_3_bits_ctrl_rfDest,
  input  [63:0] io__in_3_bits_data_src1,
  input  [63:0] io__in_3_bits_data_src2,
  input  [63:0] io__in_3_bits_data_src3,
  input  [4:0]  io__in_3_bits_InstNo,
  input         io__in_3_bits_InstFlag,
  output        io__in_4_ready,
  input         io__in_4_valid,
  input  [63:0] io__in_4_bits_cf_instr,
  input  [38:0] io__in_4_bits_cf_pc,
  input         io__in_4_bits_cf_exceptionVec_1,
  input         io__in_4_bits_cf_exceptionVec_2,
  input         io__in_4_bits_cf_exceptionVec_12,
  input         io__in_4_bits_cf_intrVec_0,
  input         io__in_4_bits_cf_intrVec_1,
  input         io__in_4_bits_cf_intrVec_2,
  input         io__in_4_bits_cf_intrVec_3,
  input         io__in_4_bits_cf_intrVec_4,
  input         io__in_4_bits_cf_intrVec_5,
  input         io__in_4_bits_cf_intrVec_6,
  input         io__in_4_bits_cf_intrVec_7,
  input         io__in_4_bits_cf_intrVec_8,
  input         io__in_4_bits_cf_intrVec_9,
  input         io__in_4_bits_cf_intrVec_10,
  input         io__in_4_bits_cf_intrVec_11,
  input         io__in_4_bits_cf_crossPageIPFFix,
  input  [63:0] io__in_4_bits_cf_runahead_checkpoint_id,
  input  [6:0]  io__in_4_bits_ctrl_fuOpType,
  input         io__in_4_bits_ctrl_rfWen,
  input  [4:0]  io__in_4_bits_ctrl_rfDest,
  input         io__in_4_bits_ctrl_isMou,
  input  [63:0] io__in_4_bits_data_src1,
  input  [63:0] io__in_4_bits_data_src2,
  input  [63:0] io__in_4_bits_data_imm,
  input  [4:0]  io__in_4_bits_InstNo,
  input         io__in_4_bits_InstFlag,
  output        io__in_5_ready,
  input         io__in_5_valid,
  input  [38:0] io__in_5_bits_cf_pc,
  input  [63:0] io__in_5_bits_cf_runahead_checkpoint_id,
  input  [6:0]  io__in_5_bits_ctrl_fuOpType,
  input         io__in_5_bits_ctrl_rfWen,
  input  [4:0]  io__in_5_bits_ctrl_rfDest,
  input  [63:0] io__in_5_bits_data_src1,
  input  [63:0] io__in_5_bits_data_src2,
  input  [4:0]  io__in_5_bits_InstNo,
  output        io__in_6_ready,
  input         io__in_6_valid,
  input  [63:0] io__in_6_bits_cf_instr,
  input  [38:0] io__in_6_bits_cf_pc,
  input  [38:0] io__in_6_bits_cf_pnpc,
  input  [3:0]  io__in_6_bits_cf_brIdx,
  input  [63:0] io__in_6_bits_cf_runahead_checkpoint_id,
  input  [6:0]  io__in_6_bits_ctrl_fuOpType,
  input         io__in_6_bits_ctrl_rfWen,
  input  [4:0]  io__in_6_bits_ctrl_rfDest,
  input  [63:0] io__in_6_bits_data_src1,
  input  [63:0] io__in_6_bits_data_src2,
  input  [63:0] io__in_6_bits_data_imm,
  input  [4:0]  io__in_6_bits_InstNo,
  output        io__in_7_ready,
  input         io__in_7_valid,
  input  [63:0] io__in_7_bits_cf_instr,
  input  [38:0] io__in_7_bits_cf_pc,
  input  [38:0] io__in_7_bits_cf_pnpc,
  input  [3:0]  io__in_7_bits_cf_brIdx,
  input  [63:0] io__in_7_bits_cf_runahead_checkpoint_id,
  input  [6:0]  io__in_7_bits_ctrl_fuOpType,
  input         io__in_7_bits_ctrl_rfWen,
  input  [4:0]  io__in_7_bits_ctrl_rfDest,
  input  [63:0] io__in_7_bits_data_src1,
  input  [63:0] io__in_7_bits_data_src2,
  input  [63:0] io__in_7_bits_data_imm,
  input  [4:0]  io__in_7_bits_InstNo,
  input         io__out_0_ready,
  output        io__out_0_valid,
  output [38:0] io__out_0_bits_decode_cf_pc,
  output [38:0] io__out_0_bits_decode_cf_redirect_target,
  output        io__out_0_bits_decode_cf_redirect_valid,
  output [63:0] io__out_0_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_0_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_0_bits_decode_ctrl_rfDest,
  output [4:0]  io__out_0_bits_decode_InstNo,
  output        io__out_0_bits_decode_InstFlag,
  output [63:0] io__out_0_bits_commits,
  input         io__out_1_ready,
  output        io__out_1_valid,
  output [38:0] io__out_1_bits_decode_cf_pc,
  output [38:0] io__out_1_bits_decode_cf_redirect_target,
  output        io__out_1_bits_decode_cf_redirect_valid,
  output [63:0] io__out_1_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_1_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_1_bits_decode_ctrl_rfDest,
  output [4:0]  io__out_1_bits_decode_InstNo,
  output        io__out_1_bits_decode_InstFlag,
  output [63:0] io__out_1_bits_commits,
  input         io__out_2_ready,
  output        io__out_2_valid,
  output [38:0] io__out_2_bits_decode_cf_pc,
  output [63:0] io__out_2_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_2_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_2_bits_decode_ctrl_rfDest,
  output        io__out_2_bits_decode_pext_OV,
  output [4:0]  io__out_2_bits_decode_InstNo,
  output [63:0] io__out_2_bits_commits,
  input         io__out_3_ready,
  output        io__out_3_valid,
  output [38:0] io__out_3_bits_decode_cf_pc,
  output [63:0] io__out_3_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_3_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_3_bits_decode_ctrl_rfDest,
  output        io__out_3_bits_decode_pext_OV,
  output [4:0]  io__out_3_bits_decode_InstNo,
  output [63:0] io__out_3_bits_commits,
  input         io__out_4_ready,
  output        io__out_4_valid,
  output [38:0] io__out_4_bits_decode_cf_pc,
  output [63:0] io__out_4_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_4_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_4_bits_decode_ctrl_rfDest,
  output [4:0]  io__out_4_bits_decode_InstNo,
  output [63:0] io__out_4_bits_commits,
  input         io__out_5_ready,
  output        io__out_5_valid,
  output [38:0] io__out_5_bits_decode_cf_pc,
  output [63:0] io__out_5_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_5_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_5_bits_decode_ctrl_rfDest,
  output [4:0]  io__out_5_bits_decode_InstNo,
  output [63:0] io__out_5_bits_commits,
  input         io__out_6_ready,
  output        io__out_6_valid,
  output [38:0] io__out_6_bits_decode_cf_pc,
  output [38:0] io__out_6_bits_decode_cf_redirect_target,
  output        io__out_6_bits_decode_cf_redirect_valid,
  output [63:0] io__out_6_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_6_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_6_bits_decode_ctrl_rfDest,
  output [4:0]  io__out_6_bits_decode_InstNo,
  output [63:0] io__out_6_bits_commits,
  input         io__out_7_ready,
  output        io__out_7_valid,
  output [38:0] io__out_7_bits_decode_cf_pc,
  output [38:0] io__out_7_bits_decode_cf_redirect_target,
  output        io__out_7_bits_decode_cf_redirect_valid,
  output [63:0] io__out_7_bits_decode_cf_runahead_checkpoint_id,
  output        io__out_7_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_7_bits_decode_ctrl_rfDest,
  output [4:0]  io__out_7_bits_decode_InstNo,
  output [63:0] io__out_7_bits_commits,
  input         io__flush,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__forward_0_valid,
  output        io__forward_0_wb_rfWen,
  output [4:0]  io__forward_0_wb_rfDest,
  output [63:0] io__forward_0_wb_rfData,
  output [4:0]  io__forward_0_InstNo,
  output        io__forward_1_valid,
  output        io__forward_1_wb_rfWen,
  output [4:0]  io__forward_1_wb_rfDest,
  output [63:0] io__forward_1_wb_rfData,
  output [4:0]  io__forward_1_InstNo,
  output        io__forward_2_valid,
  output        io__forward_2_wb_rfWen,
  output [4:0]  io__forward_2_wb_rfDest,
  output [63:0] io__forward_2_wb_rfData,
  output [4:0]  io__forward_2_InstNo,
  output        io__forward_3_valid,
  output        io__forward_3_wb_rfWen,
  output [4:0]  io__forward_3_wb_rfDest,
  output [63:0] io__forward_3_wb_rfData,
  output [4:0]  io__forward_3_InstNo,
  output        io__forward_4_valid,
  output        io__forward_4_wb_rfWen,
  output [4:0]  io__forward_4_wb_rfDest,
  output [63:0] io__forward_4_wb_rfData,
  output [4:0]  io__forward_4_InstNo,
  output        io__forward_5_valid,
  output        io__forward_5_wb_rfWen,
  output [4:0]  io__forward_5_wb_rfDest,
  output [63:0] io__forward_5_wb_rfData,
  output [4:0]  io__forward_5_InstNo,
  output        io__forward_6_valid,
  output        io__forward_6_wb_rfWen,
  output [4:0]  io__forward_6_wb_rfDest,
  output [63:0] io__forward_6_wb_rfData,
  output [4:0]  io__forward_6_InstNo,
  output        io__forward_7_valid,
  output        io__forward_7_wb_rfWen,
  output [4:0]  io__forward_7_wb_rfDest,
  output [63:0] io__forward_7_wb_rfData,
  output [4:0]  io__forward_7_InstNo,
  output [1:0]  io__memMMU_imem_priviledgeMode,
  output [1:0]  io__memMMU_dmem_priviledgeMode,
  output        io__memMMU_dmem_status_sum,
  output        io__memMMU_dmem_status_mxr,
  input         io__memMMU_dmem_loadPF,
  input         io__memMMU_dmem_storePF,
  input  [38:0] io__memMMU_dmem_addr,
  output        lsu_firststage_fire,
  input         _T_408,
  input         _T_137_0,
  output        flushICache,
  input         _T_140_0,
  output [63:0] perfCnts_2,
  output        _WIRE_2_0,
  output [63:0] satp,
  output        bpuUpdateReq_valid,
  output [38:0] bpuUpdateReq_pc,
  output        bpuUpdateReq_isMissPredict,
  output [38:0] bpuUpdateReq_actualTarget,
  output        bpuUpdateReq_actualTaken,
  output [6:0]  bpuUpdateReq_fuOpType,
  output [1:0]  bpuUpdateReq_btbType,
  output        bpuUpdateReq_isRVC,
  input         io_in_0_valid,
  input         ismmio,
  input         _WIRE_2_1,
  input         io_extra_mtip,
  output        amoReq,
  input         _T_136_0,
  input         io_extra_meip_0,
  input         _T_139_0,
  input         vmEnable,
  output [63:0] intrVec,
  input         _T_407,
  output        _WIRE_1_0,
  input         io_extra_msip,
  input         _T_138_0,
  output        flushTLB,
  input         _T_135_0
);
  wire  alu_clock; // @[SIMD_EXU.scala 212:19]
  wire  alu_reset; // @[SIMD_EXU.scala 212:19]
  wire  alu_io_in_valid; // @[SIMD_EXU.scala 212:19]
  wire [63:0] alu_io_in_bits_src1; // @[SIMD_EXU.scala 212:19]
  wire [63:0] alu_io_in_bits_src2; // @[SIMD_EXU.scala 212:19]
  wire [6:0] alu_io_in_bits_func; // @[SIMD_EXU.scala 212:19]
  wire [63:0] alu_io_out_bits; // @[SIMD_EXU.scala 212:19]
  wire [63:0] alu_io_cfIn_instr; // @[SIMD_EXU.scala 212:19]
  wire [38:0] alu_io_cfIn_pc; // @[SIMD_EXU.scala 212:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[SIMD_EXU.scala 212:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[SIMD_EXU.scala 212:19]
  wire [38:0] alu_io_redirect_target; // @[SIMD_EXU.scala 212:19]
  wire  alu_io_redirect_valid; // @[SIMD_EXU.scala 212:19]
  wire [63:0] alu_io_offset; // @[SIMD_EXU.scala 212:19]
  wire  alu1_clock; // @[SIMD_EXU.scala 222:20]
  wire  alu1_reset; // @[SIMD_EXU.scala 222:20]
  wire  alu1_io_in_valid; // @[SIMD_EXU.scala 222:20]
  wire [63:0] alu1_io_in_bits_src1; // @[SIMD_EXU.scala 222:20]
  wire [63:0] alu1_io_in_bits_src2; // @[SIMD_EXU.scala 222:20]
  wire [6:0] alu1_io_in_bits_func; // @[SIMD_EXU.scala 222:20]
  wire [63:0] alu1_io_out_bits; // @[SIMD_EXU.scala 222:20]
  wire [63:0] alu1_io_cfIn_instr; // @[SIMD_EXU.scala 222:20]
  wire [38:0] alu1_io_cfIn_pc; // @[SIMD_EXU.scala 222:20]
  wire [38:0] alu1_io_cfIn_pnpc; // @[SIMD_EXU.scala 222:20]
  wire [3:0] alu1_io_cfIn_brIdx; // @[SIMD_EXU.scala 222:20]
  wire [38:0] alu1_io_redirect_target; // @[SIMD_EXU.scala 222:20]
  wire  alu1_io_redirect_valid; // @[SIMD_EXU.scala 222:20]
  wire [63:0] alu1_io_offset; // @[SIMD_EXU.scala 222:20]
  wire  SIMDU_2way_clock; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_reset; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_flush; // @[SIMD_EXU.scala 232:23]
  wire [38:0] SIMDU_2way_io_DecodeOut_0_cf_pc; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeOut_0_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeOut_0_ctrl_rfWen; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeOut_0_ctrl_rfDest; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeOut_0_pext_OV; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeOut_0_InstNo; // @[SIMD_EXU.scala 232:23]
  wire [38:0] SIMDU_2way_io_DecodeOut_1_cf_pc; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeOut_1_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeOut_1_ctrl_rfWen; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeOut_1_ctrl_rfDest; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeOut_1_pext_OV; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeOut_1_InstNo; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_0_cf_instr; // @[SIMD_EXU.scala 232:23]
  wire [38:0] SIMDU_2way_io_DecodeIn_0_cf_pc; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_0_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeIn_0_cf_instrType; // @[SIMD_EXU.scala 232:23]
  wire [6:0] SIMDU_2way_io_DecodeIn_0_ctrl_fuOpType; // @[SIMD_EXU.scala 232:23]
  wire [2:0] SIMDU_2way_io_DecodeIn_0_ctrl_funct3; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_0_ctrl_func24; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_0_ctrl_func23; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_0_ctrl_rfWen; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeIn_0_ctrl_rfDest; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_0_data_src1; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_0_data_src2; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_0_data_src3; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeIn_0_InstNo; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_0_InstFlag; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_1_cf_instr; // @[SIMD_EXU.scala 232:23]
  wire [38:0] SIMDU_2way_io_DecodeIn_1_cf_pc; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_1_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeIn_1_cf_instrType; // @[SIMD_EXU.scala 232:23]
  wire [6:0] SIMDU_2way_io_DecodeIn_1_ctrl_fuOpType; // @[SIMD_EXU.scala 232:23]
  wire [2:0] SIMDU_2way_io_DecodeIn_1_ctrl_funct3; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_1_ctrl_func24; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_1_ctrl_func23; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_1_ctrl_rfWen; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeIn_1_ctrl_rfDest; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_1_data_src1; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_1_data_src2; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_DecodeIn_1_data_src3; // @[SIMD_EXU.scala 232:23]
  wire [4:0] SIMDU_2way_io_DecodeIn_1_InstNo; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_DecodeIn_1_InstFlag; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_FirstStageFire_0; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_FirstStageFire_1; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_in_0_ready; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_in_0_valid; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_in_1_ready; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_in_1_valid; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_out_0_ready; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_out_0_valid; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_out_0_bits; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_out_1_ready; // @[SIMD_EXU.scala 232:23]
  wire  SIMDU_2way_io_out_1_valid; // @[SIMD_EXU.scala 232:23]
  wire [63:0] SIMDU_2way_io_out_1_bits; // @[SIMD_EXU.scala 232:23]
  wire  mdu_clock; // @[SIMD_EXU.scala 277:19]
  wire  mdu_reset; // @[SIMD_EXU.scala 277:19]
  wire  mdu_io_in_ready; // @[SIMD_EXU.scala 277:19]
  wire  mdu_io_in_valid; // @[SIMD_EXU.scala 277:19]
  wire [63:0] mdu_io_in_bits_src1; // @[SIMD_EXU.scala 277:19]
  wire [63:0] mdu_io_in_bits_src2; // @[SIMD_EXU.scala 277:19]
  wire [6:0] mdu_io_in_bits_func; // @[SIMD_EXU.scala 277:19]
  wire  mdu_io_out_ready; // @[SIMD_EXU.scala 277:19]
  wire  mdu_io_out_valid; // @[SIMD_EXU.scala 277:19]
  wire [63:0] mdu_io_out_bits; // @[SIMD_EXU.scala 277:19]
  wire  mdu_io_flush; // @[SIMD_EXU.scala 277:19]
  wire  ALU_clock; // @[SIMD_EXU.scala 285:21]
  wire  ALU_reset; // @[SIMD_EXU.scala 285:21]
  wire  ALU_io_in_valid; // @[SIMD_EXU.scala 285:21]
  wire [63:0] ALU_io_in_bits_src1; // @[SIMD_EXU.scala 285:21]
  wire [63:0] ALU_io_in_bits_src2; // @[SIMD_EXU.scala 285:21]
  wire [6:0] ALU_io_in_bits_func; // @[SIMD_EXU.scala 285:21]
  wire  ALU_io_out_ready; // @[SIMD_EXU.scala 285:21]
  wire  ALU_io_out_valid; // @[SIMD_EXU.scala 285:21]
  wire [63:0] ALU_io_out_bits; // @[SIMD_EXU.scala 285:21]
  wire [63:0] ALU_io_cfIn_instr; // @[SIMD_EXU.scala 285:21]
  wire [38:0] ALU_io_cfIn_pc; // @[SIMD_EXU.scala 285:21]
  wire [38:0] ALU_io_cfIn_pnpc; // @[SIMD_EXU.scala 285:21]
  wire [3:0] ALU_io_cfIn_brIdx; // @[SIMD_EXU.scala 285:21]
  wire [38:0] ALU_io_redirect_target; // @[SIMD_EXU.scala 285:21]
  wire  ALU_io_redirect_valid; // @[SIMD_EXU.scala 285:21]
  wire [63:0] ALU_io_offset; // @[SIMD_EXU.scala 285:21]
  wire  ALU_bpuUpdateReq_0_valid; // @[SIMD_EXU.scala 285:21]
  wire [38:0] ALU_bpuUpdateReq_0_pc; // @[SIMD_EXU.scala 285:21]
  wire  ALU_bpuUpdateReq_0_isMissPredict; // @[SIMD_EXU.scala 285:21]
  wire [38:0] ALU_bpuUpdateReq_0_actualTarget; // @[SIMD_EXU.scala 285:21]
  wire  ALU_bpuUpdateReq_0_actualTaken; // @[SIMD_EXU.scala 285:21]
  wire [6:0] ALU_bpuUpdateReq_0_fuOpType; // @[SIMD_EXU.scala 285:21]
  wire [1:0] ALU_bpuUpdateReq_0_btbType; // @[SIMD_EXU.scala 285:21]
  wire  ALU_bpuUpdateReq_0_isRVC; // @[SIMD_EXU.scala 285:21]
  wire  lsu_clock; // @[SIMD_EXU.scala 298:19]
  wire  lsu_reset; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_in_ready; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_in_valid; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_in_bits_src1; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_in_bits_src2; // @[SIMD_EXU.scala 298:19]
  wire [6:0] lsu_io_in_bits_func; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_out_ready; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_out_valid; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_out_bits; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_wdata; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_dmem_req_ready; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_dmem_req_valid; // @[SIMD_EXU.scala 298:19]
  wire [38:0] lsu_io_dmem_req_bits_addr; // @[SIMD_EXU.scala 298:19]
  wire [2:0] lsu_io_dmem_req_bits_size; // @[SIMD_EXU.scala 298:19]
  wire [3:0] lsu_io_dmem_req_bits_cmd; // @[SIMD_EXU.scala 298:19]
  wire [7:0] lsu_io_dmem_req_bits_wmask; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_dmem_req_bits_wdata; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_dmem_resp_valid; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_dmem_resp_bits_rdata; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_loadAddrMisaligned; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_storeAddrMisaligned; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_flush; // @[SIMD_EXU.scala 298:19]
  wire [38:0] lsu_io_DecodeOut_cf_pc; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_exceptionVec_1; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_exceptionVec_2; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_exceptionVec_12; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_0; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_1; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_2; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_3; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_4; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_5; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_6; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_7; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_8; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_9; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_10; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_intrVec_11; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_cf_crossPageIPFFix; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_DecodeOut_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_ctrl_rfWen; // @[SIMD_EXU.scala 298:19]
  wire [4:0] lsu_io_DecodeOut_ctrl_rfDest; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_ctrl_isMou; // @[SIMD_EXU.scala 298:19]
  wire [4:0] lsu_io_DecodeOut_InstNo; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeOut_InstFlag; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_DecodeIn_cf_instr; // @[SIMD_EXU.scala 298:19]
  wire [38:0] lsu_io_DecodeIn_cf_pc; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_exceptionVec_1; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_exceptionVec_2; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_exceptionVec_12; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_0; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_1; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_2; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_3; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_4; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_5; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_6; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_7; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_8; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_9; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_10; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_intrVec_11; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_cf_crossPageIPFFix; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_io_DecodeIn_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_ctrl_rfWen; // @[SIMD_EXU.scala 298:19]
  wire [4:0] lsu_io_DecodeIn_ctrl_rfDest; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_ctrl_isMou; // @[SIMD_EXU.scala 298:19]
  wire [4:0] lsu_io_DecodeIn_InstNo; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_DecodeIn_InstFlag; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_loadPF; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_storePF; // @[SIMD_EXU.scala 298:19]
  wire  lsu_lsu_firststage_fire_0; // @[SIMD_EXU.scala 298:19]
  wire  lsu_setLr; // @[SIMD_EXU.scala 298:19]
  wire  lsu__T_408; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_memMMU_dmem_loadPF; // @[SIMD_EXU.scala 298:19]
  wire  lsu_ismmio; // @[SIMD_EXU.scala 298:19]
  wire  lsu_lr; // @[SIMD_EXU.scala 298:19]
  wire  lsu_amoReq; // @[SIMD_EXU.scala 298:19]
  wire  lsu_io_memMMU_dmem_storePF; // @[SIMD_EXU.scala 298:19]
  wire  lsu_vmEnable; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_addr_0; // @[SIMD_EXU.scala 298:19]
  wire  lsu__T_407; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_setLrAddr; // @[SIMD_EXU.scala 298:19]
  wire  lsu_setLrVal; // @[SIMD_EXU.scala 298:19]
  wire [63:0] lsu_lrAddr; // @[SIMD_EXU.scala 298:19]
  wire  csr_clock; // @[SIMD_EXU.scala 315:19]
  wire  csr_reset; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_in_valid; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_io_in_bits_src1; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_io_in_bits_src2; // @[SIMD_EXU.scala 315:19]
  wire [6:0] csr_io_in_bits_func; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_io_out_bits; // @[SIMD_EXU.scala 315:19]
  wire [38:0] csr_io_cfIn_pc; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_13; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_exceptionVec_15; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_0; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_1; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_2; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_3; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_4; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_5; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_6; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_7; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_8; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_9; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_10; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_intrVec_11; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_cfIn_crossPageIPFFix; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_ctrlIn_isMou; // @[SIMD_EXU.scala 315:19]
  wire [38:0] csr_io_redirect_target; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_redirect_valid; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_instrValid; // @[SIMD_EXU.scala 315:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[SIMD_EXU.scala 315:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_dmemMMU_status_sum; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_dmemMMU_status_mxr; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_dmemMMU_loadPF; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_dmemMMU_storePF; // @[SIMD_EXU.scala 315:19]
  wire [38:0] csr_io_dmemMMU_addr; // @[SIMD_EXU.scala 315:19]
  wire  csr_io_wenFix; // @[SIMD_EXU.scala 315:19]
  wire  csr_set_lr; // @[SIMD_EXU.scala 315:19]
  wire  csr_flushICache_0; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_satp_0; // @[SIMD_EXU.scala 315:19]
  wire  csr_lr_0; // @[SIMD_EXU.scala 315:19]
  wire  csr_OVWEN_0; // @[SIMD_EXU.scala 315:19]
  wire  csr_mtip; // @[SIMD_EXU.scala 315:19]
  wire  csr_meip; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_LSUADDR; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_intrVec_0; // @[SIMD_EXU.scala 315:19]
  wire  csr_msip; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_set_lr_addr; // @[SIMD_EXU.scala 315:19]
  wire  csr_flushTLB_0; // @[SIMD_EXU.scala 315:19]
  wire  csr_set_lr_val; // @[SIMD_EXU.scala 315:19]
  wire [63:0] csr_lrAddr_0; // @[SIMD_EXU.scala 315:19]
  wire  PerfU_clock; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_reset; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMultiCommit3; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMultiCommit6; // @[SIMD_EXU.scala 362:21]
  wire [63:0] PerfU_perfCnts_2_0; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMinstret; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMultiCommit2; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMultiCommit5; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMultiCommit4; // @[SIMD_EXU.scala 362:21]
  wire  PerfU_perfCntCondMultiCommit; // @[SIMD_EXU.scala 362:21]
  wire  _T_1 = io__out_0_ready & io__out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io__out_1_ready & io__out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_16 = io__out_5_ready & io__out_5_valid; // @[Decoupled.scala 40:37]
  wire  _T_19 = io__out_6_ready & io__out_6_valid; // @[Decoupled.scala 40:37]
  wire  _T_22 = io__out_7_ready & io__out_7_valid; // @[Decoupled.scala 40:37]
  wire  _T_37 = io__in_0_bits_InstNo <= io__in_4_bits_InstNo & io__in_0_bits_InstFlag == io__in_4_bits_InstFlag |
    io__in_0_bits_InstNo > io__in_4_bits_InstNo & io__in_0_bits_InstFlag != io__in_4_bits_InstFlag; // @[SIMD_EXU.scala 188:101]
  wire  BeforeLSUhasRedirect = _T_37 & io__out_0_bits_decode_cf_redirect_valid; // @[SIMD_EXU.scala 297:147]
  wire [38:0] csr_bits_cf_pc = io__in_1_valid ? io__in_1_bits_cf_pc : lsu_io_DecodeOut_cf_pc; // @[SIMD_EXU.scala 314:21]
  wire [63:0] csr_bits_cf_runahead_checkpoint_id = io__in_1_valid ? io__in_1_bits_cf_runahead_checkpoint_id :
    lsu_io_DecodeOut_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 314:21]
  wire  csr_bits_ctrl_rfWen = io__in_1_valid ? io__in_1_bits_ctrl_rfWen : lsu_io_DecodeOut_ctrl_rfWen; // @[SIMD_EXU.scala 314:21]
  wire [4:0] csr_bits_ctrl_rfDest = io__in_1_valid ? io__in_1_bits_ctrl_rfDest : lsu_io_DecodeOut_ctrl_rfDest; // @[SIMD_EXU.scala 314:21]
  wire [4:0] csr_bits_InstNo = io__in_1_valid ? io__in_1_bits_InstNo : lsu_io_DecodeOut_InstNo; // @[SIMD_EXU.scala 314:21]
  wire  csr_bits_InstFlag = io__in_1_valid ? io__in_1_bits_InstFlag : lsu_io_DecodeOut_InstFlag; // @[SIMD_EXU.scala 314:21]
  wire  lsuexp = lsu_io_loadAddrMisaligned | lsu_io_storeAddrMisaligned | lsu_io_storePF | lsu_io_loadPF; // @[SIMD_EXU.scala 340:87]
  wire  csrfix = csr_io_wenFix & io__in_1_valid; // @[SIMD_EXU.scala 341:31]
  wire  _GEN_15 = lsuexp ? csr_bits_ctrl_rfWen : io__in_1_bits_ctrl_rfWen; // @[SIMD_EXU.scala 352:15 355:32 203:38]
  wire  _WIRE_1 = SIMDU_2way_io_FirstStageFire_0; // @[SIMD_EXU.scala 240:37 241:27]
  wire  _WIRE_2 = SIMDU_2way_io_FirstStageFire_1; // @[SIMD_EXU.scala 243:38 244:28]
  ALU alu ( // @[SIMD_EXU.scala 212:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset)
  );
  ALU_1 alu1 ( // @[SIMD_EXU.scala 222:20]
    .clock(alu1_clock),
    .reset(alu1_reset),
    .io_in_valid(alu1_io_in_valid),
    .io_in_bits_src1(alu1_io_in_bits_src1),
    .io_in_bits_src2(alu1_io_in_bits_src2),
    .io_in_bits_func(alu1_io_in_bits_func),
    .io_out_bits(alu1_io_out_bits),
    .io_cfIn_instr(alu1_io_cfIn_instr),
    .io_cfIn_pc(alu1_io_cfIn_pc),
    .io_cfIn_pnpc(alu1_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu1_io_cfIn_brIdx),
    .io_redirect_target(alu1_io_redirect_target),
    .io_redirect_valid(alu1_io_redirect_valid),
    .io_offset(alu1_io_offset)
  );
  SIMDU_2way SIMDU_2way ( // @[SIMD_EXU.scala 232:23]
    .clock(SIMDU_2way_clock),
    .reset(SIMDU_2way_reset),
    .io_flush(SIMDU_2way_io_flush),
    .io_DecodeOut_0_cf_pc(SIMDU_2way_io_DecodeOut_0_cf_pc),
    .io_DecodeOut_0_cf_runahead_checkpoint_id(SIMDU_2way_io_DecodeOut_0_cf_runahead_checkpoint_id),
    .io_DecodeOut_0_ctrl_rfWen(SIMDU_2way_io_DecodeOut_0_ctrl_rfWen),
    .io_DecodeOut_0_ctrl_rfDest(SIMDU_2way_io_DecodeOut_0_ctrl_rfDest),
    .io_DecodeOut_0_pext_OV(SIMDU_2way_io_DecodeOut_0_pext_OV),
    .io_DecodeOut_0_InstNo(SIMDU_2way_io_DecodeOut_0_InstNo),
    .io_DecodeOut_1_cf_pc(SIMDU_2way_io_DecodeOut_1_cf_pc),
    .io_DecodeOut_1_cf_runahead_checkpoint_id(SIMDU_2way_io_DecodeOut_1_cf_runahead_checkpoint_id),
    .io_DecodeOut_1_ctrl_rfWen(SIMDU_2way_io_DecodeOut_1_ctrl_rfWen),
    .io_DecodeOut_1_ctrl_rfDest(SIMDU_2way_io_DecodeOut_1_ctrl_rfDest),
    .io_DecodeOut_1_pext_OV(SIMDU_2way_io_DecodeOut_1_pext_OV),
    .io_DecodeOut_1_InstNo(SIMDU_2way_io_DecodeOut_1_InstNo),
    .io_DecodeIn_0_cf_instr(SIMDU_2way_io_DecodeIn_0_cf_instr),
    .io_DecodeIn_0_cf_pc(SIMDU_2way_io_DecodeIn_0_cf_pc),
    .io_DecodeIn_0_cf_runahead_checkpoint_id(SIMDU_2way_io_DecodeIn_0_cf_runahead_checkpoint_id),
    .io_DecodeIn_0_cf_instrType(SIMDU_2way_io_DecodeIn_0_cf_instrType),
    .io_DecodeIn_0_ctrl_fuOpType(SIMDU_2way_io_DecodeIn_0_ctrl_fuOpType),
    .io_DecodeIn_0_ctrl_funct3(SIMDU_2way_io_DecodeIn_0_ctrl_funct3),
    .io_DecodeIn_0_ctrl_func24(SIMDU_2way_io_DecodeIn_0_ctrl_func24),
    .io_DecodeIn_0_ctrl_func23(SIMDU_2way_io_DecodeIn_0_ctrl_func23),
    .io_DecodeIn_0_ctrl_rfWen(SIMDU_2way_io_DecodeIn_0_ctrl_rfWen),
    .io_DecodeIn_0_ctrl_rfDest(SIMDU_2way_io_DecodeIn_0_ctrl_rfDest),
    .io_DecodeIn_0_data_src1(SIMDU_2way_io_DecodeIn_0_data_src1),
    .io_DecodeIn_0_data_src2(SIMDU_2way_io_DecodeIn_0_data_src2),
    .io_DecodeIn_0_data_src3(SIMDU_2way_io_DecodeIn_0_data_src3),
    .io_DecodeIn_0_InstNo(SIMDU_2way_io_DecodeIn_0_InstNo),
    .io_DecodeIn_0_InstFlag(SIMDU_2way_io_DecodeIn_0_InstFlag),
    .io_DecodeIn_1_cf_instr(SIMDU_2way_io_DecodeIn_1_cf_instr),
    .io_DecodeIn_1_cf_pc(SIMDU_2way_io_DecodeIn_1_cf_pc),
    .io_DecodeIn_1_cf_runahead_checkpoint_id(SIMDU_2way_io_DecodeIn_1_cf_runahead_checkpoint_id),
    .io_DecodeIn_1_cf_instrType(SIMDU_2way_io_DecodeIn_1_cf_instrType),
    .io_DecodeIn_1_ctrl_fuOpType(SIMDU_2way_io_DecodeIn_1_ctrl_fuOpType),
    .io_DecodeIn_1_ctrl_funct3(SIMDU_2way_io_DecodeIn_1_ctrl_funct3),
    .io_DecodeIn_1_ctrl_func24(SIMDU_2way_io_DecodeIn_1_ctrl_func24),
    .io_DecodeIn_1_ctrl_func23(SIMDU_2way_io_DecodeIn_1_ctrl_func23),
    .io_DecodeIn_1_ctrl_rfWen(SIMDU_2way_io_DecodeIn_1_ctrl_rfWen),
    .io_DecodeIn_1_ctrl_rfDest(SIMDU_2way_io_DecodeIn_1_ctrl_rfDest),
    .io_DecodeIn_1_data_src1(SIMDU_2way_io_DecodeIn_1_data_src1),
    .io_DecodeIn_1_data_src2(SIMDU_2way_io_DecodeIn_1_data_src2),
    .io_DecodeIn_1_data_src3(SIMDU_2way_io_DecodeIn_1_data_src3),
    .io_DecodeIn_1_InstNo(SIMDU_2way_io_DecodeIn_1_InstNo),
    .io_DecodeIn_1_InstFlag(SIMDU_2way_io_DecodeIn_1_InstFlag),
    .io_FirstStageFire_0(SIMDU_2way_io_FirstStageFire_0),
    .io_FirstStageFire_1(SIMDU_2way_io_FirstStageFire_1),
    .io_in_0_ready(SIMDU_2way_io_in_0_ready),
    .io_in_0_valid(SIMDU_2way_io_in_0_valid),
    .io_in_1_ready(SIMDU_2way_io_in_1_ready),
    .io_in_1_valid(SIMDU_2way_io_in_1_valid),
    .io_out_0_ready(SIMDU_2way_io_out_0_ready),
    .io_out_0_valid(SIMDU_2way_io_out_0_valid),
    .io_out_0_bits(SIMDU_2way_io_out_0_bits),
    .io_out_1_ready(SIMDU_2way_io_out_1_ready),
    .io_out_1_valid(SIMDU_2way_io_out_1_valid),
    .io_out_1_bits(SIMDU_2way_io_out_1_bits)
  );
  MDU mdu ( // @[SIMD_EXU.scala 277:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits),
    .io_flush(mdu_io_flush)
  );
  ALU_2 ALU ( // @[SIMD_EXU.scala 285:21]
    .clock(ALU_clock),
    .reset(ALU_reset),
    .io_in_valid(ALU_io_in_valid),
    .io_in_bits_src1(ALU_io_in_bits_src1),
    .io_in_bits_src2(ALU_io_in_bits_src2),
    .io_in_bits_func(ALU_io_in_bits_func),
    .io_out_ready(ALU_io_out_ready),
    .io_out_valid(ALU_io_out_valid),
    .io_out_bits(ALU_io_out_bits),
    .io_cfIn_instr(ALU_io_cfIn_instr),
    .io_cfIn_pc(ALU_io_cfIn_pc),
    .io_cfIn_pnpc(ALU_io_cfIn_pnpc),
    .io_cfIn_brIdx(ALU_io_cfIn_brIdx),
    .io_redirect_target(ALU_io_redirect_target),
    .io_redirect_valid(ALU_io_redirect_valid),
    .io_offset(ALU_io_offset),
    .bpuUpdateReq_0_valid(ALU_bpuUpdateReq_0_valid),
    .bpuUpdateReq_0_pc(ALU_bpuUpdateReq_0_pc),
    .bpuUpdateReq_0_isMissPredict(ALU_bpuUpdateReq_0_isMissPredict),
    .bpuUpdateReq_0_actualTarget(ALU_bpuUpdateReq_0_actualTarget),
    .bpuUpdateReq_0_actualTaken(ALU_bpuUpdateReq_0_actualTaken),
    .bpuUpdateReq_0_fuOpType(ALU_bpuUpdateReq_0_fuOpType),
    .bpuUpdateReq_0_btbType(ALU_bpuUpdateReq_0_btbType),
    .bpuUpdateReq_0_isRVC(ALU_bpuUpdateReq_0_isRVC)
  );
  pipeline_lsu_atom lsu ( // @[SIMD_EXU.scala 298:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_in_ready(lsu_io_in_ready),
    .io_in_valid(lsu_io_in_valid),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .io_in_bits_src2(lsu_io_in_bits_src2),
    .io_in_bits_func(lsu_io_in_bits_func),
    .io_out_ready(lsu_io_out_ready),
    .io_out_valid(lsu_io_out_valid),
    .io_out_bits(lsu_io_out_bits),
    .io_wdata(lsu_io_wdata),
    .io_dmem_req_ready(lsu_io_dmem_req_ready),
    .io_dmem_req_valid(lsu_io_dmem_req_valid),
    .io_dmem_req_bits_addr(lsu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(lsu_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(lsu_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(lsu_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(lsu_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(lsu_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(lsu_io_dmem_resp_bits_rdata),
    .io_loadAddrMisaligned(lsu_io_loadAddrMisaligned),
    .io_storeAddrMisaligned(lsu_io_storeAddrMisaligned),
    .io_flush(lsu_io_flush),
    .io_DecodeOut_cf_pc(lsu_io_DecodeOut_cf_pc),
    .io_DecodeOut_cf_exceptionVec_1(lsu_io_DecodeOut_cf_exceptionVec_1),
    .io_DecodeOut_cf_exceptionVec_2(lsu_io_DecodeOut_cf_exceptionVec_2),
    .io_DecodeOut_cf_exceptionVec_12(lsu_io_DecodeOut_cf_exceptionVec_12),
    .io_DecodeOut_cf_intrVec_0(lsu_io_DecodeOut_cf_intrVec_0),
    .io_DecodeOut_cf_intrVec_1(lsu_io_DecodeOut_cf_intrVec_1),
    .io_DecodeOut_cf_intrVec_2(lsu_io_DecodeOut_cf_intrVec_2),
    .io_DecodeOut_cf_intrVec_3(lsu_io_DecodeOut_cf_intrVec_3),
    .io_DecodeOut_cf_intrVec_4(lsu_io_DecodeOut_cf_intrVec_4),
    .io_DecodeOut_cf_intrVec_5(lsu_io_DecodeOut_cf_intrVec_5),
    .io_DecodeOut_cf_intrVec_6(lsu_io_DecodeOut_cf_intrVec_6),
    .io_DecodeOut_cf_intrVec_7(lsu_io_DecodeOut_cf_intrVec_7),
    .io_DecodeOut_cf_intrVec_8(lsu_io_DecodeOut_cf_intrVec_8),
    .io_DecodeOut_cf_intrVec_9(lsu_io_DecodeOut_cf_intrVec_9),
    .io_DecodeOut_cf_intrVec_10(lsu_io_DecodeOut_cf_intrVec_10),
    .io_DecodeOut_cf_intrVec_11(lsu_io_DecodeOut_cf_intrVec_11),
    .io_DecodeOut_cf_crossPageIPFFix(lsu_io_DecodeOut_cf_crossPageIPFFix),
    .io_DecodeOut_cf_runahead_checkpoint_id(lsu_io_DecodeOut_cf_runahead_checkpoint_id),
    .io_DecodeOut_ctrl_rfWen(lsu_io_DecodeOut_ctrl_rfWen),
    .io_DecodeOut_ctrl_rfDest(lsu_io_DecodeOut_ctrl_rfDest),
    .io_DecodeOut_ctrl_isMou(lsu_io_DecodeOut_ctrl_isMou),
    .io_DecodeOut_InstNo(lsu_io_DecodeOut_InstNo),
    .io_DecodeOut_InstFlag(lsu_io_DecodeOut_InstFlag),
    .io_DecodeIn_cf_instr(lsu_io_DecodeIn_cf_instr),
    .io_DecodeIn_cf_pc(lsu_io_DecodeIn_cf_pc),
    .io_DecodeIn_cf_exceptionVec_1(lsu_io_DecodeIn_cf_exceptionVec_1),
    .io_DecodeIn_cf_exceptionVec_2(lsu_io_DecodeIn_cf_exceptionVec_2),
    .io_DecodeIn_cf_exceptionVec_12(lsu_io_DecodeIn_cf_exceptionVec_12),
    .io_DecodeIn_cf_intrVec_0(lsu_io_DecodeIn_cf_intrVec_0),
    .io_DecodeIn_cf_intrVec_1(lsu_io_DecodeIn_cf_intrVec_1),
    .io_DecodeIn_cf_intrVec_2(lsu_io_DecodeIn_cf_intrVec_2),
    .io_DecodeIn_cf_intrVec_3(lsu_io_DecodeIn_cf_intrVec_3),
    .io_DecodeIn_cf_intrVec_4(lsu_io_DecodeIn_cf_intrVec_4),
    .io_DecodeIn_cf_intrVec_5(lsu_io_DecodeIn_cf_intrVec_5),
    .io_DecodeIn_cf_intrVec_6(lsu_io_DecodeIn_cf_intrVec_6),
    .io_DecodeIn_cf_intrVec_7(lsu_io_DecodeIn_cf_intrVec_7),
    .io_DecodeIn_cf_intrVec_8(lsu_io_DecodeIn_cf_intrVec_8),
    .io_DecodeIn_cf_intrVec_9(lsu_io_DecodeIn_cf_intrVec_9),
    .io_DecodeIn_cf_intrVec_10(lsu_io_DecodeIn_cf_intrVec_10),
    .io_DecodeIn_cf_intrVec_11(lsu_io_DecodeIn_cf_intrVec_11),
    .io_DecodeIn_cf_crossPageIPFFix(lsu_io_DecodeIn_cf_crossPageIPFFix),
    .io_DecodeIn_cf_runahead_checkpoint_id(lsu_io_DecodeIn_cf_runahead_checkpoint_id),
    .io_DecodeIn_ctrl_rfWen(lsu_io_DecodeIn_ctrl_rfWen),
    .io_DecodeIn_ctrl_rfDest(lsu_io_DecodeIn_ctrl_rfDest),
    .io_DecodeIn_ctrl_isMou(lsu_io_DecodeIn_ctrl_isMou),
    .io_DecodeIn_InstNo(lsu_io_DecodeIn_InstNo),
    .io_DecodeIn_InstFlag(lsu_io_DecodeIn_InstFlag),
    .io_loadPF(lsu_io_loadPF),
    .io_storePF(lsu_io_storePF),
    .lsu_firststage_fire_0(lsu_lsu_firststage_fire_0),
    .setLr(lsu_setLr),
    ._T_408(lsu__T_408),
    .io_memMMU_dmem_loadPF(lsu_io_memMMU_dmem_loadPF),
    .ismmio(lsu_ismmio),
    .lr(lsu_lr),
    .amoReq(lsu_amoReq),
    .io_memMMU_dmem_storePF(lsu_io_memMMU_dmem_storePF),
    .vmEnable(lsu_vmEnable),
    .addr_0(lsu_addr_0),
    ._T_407(lsu__T_407),
    .setLrAddr(lsu_setLrAddr),
    .setLrVal(lsu_setLrVal),
    .lrAddr(lsu_lrAddr)
  );
  new_SIMD_CSR csr ( // @[SIMD_EXU.scala 315:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_exceptionVec_13(csr_io_cfIn_exceptionVec_13),
    .io_cfIn_exceptionVec_15(csr_io_cfIn_exceptionVec_15),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossPageIPFFix(csr_io_cfIn_crossPageIPFFix),
    .io_ctrlIn_isMou(csr_io_ctrlIn_isMou),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_addr(csr_io_dmemMMU_addr),
    .io_wenFix(csr_io_wenFix),
    .set_lr(csr_set_lr),
    .flushICache_0(csr_flushICache_0),
    .satp_0(csr_satp_0),
    .lr_0(csr_lr_0),
    .OVWEN_0(csr_OVWEN_0),
    .mtip(csr_mtip),
    .meip(csr_meip),
    .LSUADDR(csr_LSUADDR),
    .intrVec_0(csr_intrVec_0),
    .msip(csr_msip),
    .set_lr_addr(csr_set_lr_addr),
    .flushTLB_0(csr_flushTLB_0),
    .set_lr_val(csr_set_lr_val),
    .lrAddr_0(csr_lrAddr_0)
  );
  PerfU PerfU ( // @[SIMD_EXU.scala 362:21]
    .clock(PerfU_clock),
    .reset(PerfU_reset),
    .perfCntCondMultiCommit3(PerfU_perfCntCondMultiCommit3),
    .perfCntCondMultiCommit6(PerfU_perfCntCondMultiCommit6),
    .perfCnts_2_0(PerfU_perfCnts_2_0),
    .perfCntCondMinstret(PerfU_perfCntCondMinstret),
    .perfCntCondMultiCommit2(PerfU_perfCntCondMultiCommit2),
    .perfCntCondMultiCommit5(PerfU_perfCntCondMultiCommit5),
    .perfCntCondMultiCommit4(PerfU_perfCntCondMultiCommit4),
    .perfCntCondMultiCommit(PerfU_perfCntCondMultiCommit)
  );
  assign io__in_0_ready = ~io__in_0_valid | _T_1; // @[SIMD_EXU.scala 206:39]
  assign io__in_1_ready = ~io__in_1_valid | _T_4; // @[SIMD_EXU.scala 206:39]
  assign io__in_2_ready = SIMDU_2way_io_in_0_ready; // @[SIMD_EXU.scala 255:28]
  assign io__in_3_ready = SIMDU_2way_io_in_1_ready; // @[SIMD_EXU.scala 256:28]
  assign io__in_4_ready = lsu_io_in_ready; // @[SIMD_EXU.scala 380:23]
  assign io__in_5_ready = ~io__in_5_valid | _T_16; // @[SIMD_EXU.scala 206:39]
  assign io__in_6_ready = ~io__in_6_valid | _T_19; // @[SIMD_EXU.scala 206:39]
  assign io__in_7_ready = ~io__in_7_valid | _T_22; // @[SIMD_EXU.scala 206:39]
  assign io__out_0_valid = io__in_0_valid; // @[SIMD_EXU.scala 291:30]
  assign io__out_0_bits_decode_cf_pc = io__in_0_bits_cf_pc; // @[SIMD_EXU.scala 202:27]
  assign io__out_0_bits_decode_cf_redirect_target = ALU_io_redirect_target; // @[SIMD_EXU.scala 290:44]
  assign io__out_0_bits_decode_cf_redirect_valid = ALU_io_redirect_valid; // @[SIMD_EXU.scala 290:44]
  assign io__out_0_bits_decode_cf_runahead_checkpoint_id = io__in_0_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 202:27]
  assign io__out_0_bits_decode_ctrl_rfWen = io__in_0_bits_ctrl_rfWen; // @[SIMD_EXU.scala 203:38]
  assign io__out_0_bits_decode_ctrl_rfDest = io__in_0_bits_ctrl_rfDest; // @[SIMD_EXU.scala 202:27]
  assign io__out_0_bits_decode_InstNo = io__in_0_bits_InstNo; // @[SIMD_EXU.scala 202:27]
  assign io__out_0_bits_decode_InstFlag = io__in_0_bits_InstFlag; // @[SIMD_EXU.scala 202:27]
  assign io__out_0_bits_commits = ALU_io_out_bits; // @[SIMD_EXU.scala 292:37]
  assign io__out_1_valid = io__in_1_valid | lsuexp; // @[SIMD_EXU.scala 372:51]
  assign io__out_1_bits_decode_cf_pc = lsuexp ? csr_bits_cf_pc : io__in_1_bits_cf_pc; // @[SIMD_EXU.scala 352:15 202:27 355:32]
  assign io__out_1_bits_decode_cf_redirect_target = csr_io_redirect_target; // @[SIMD_EXU.scala 364:42]
  assign io__out_1_bits_decode_cf_redirect_valid = csr_io_redirect_valid; // @[SIMD_EXU.scala 364:42]
  assign io__out_1_bits_decode_cf_runahead_checkpoint_id = lsuexp ? csr_bits_cf_runahead_checkpoint_id :
    io__in_1_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 352:15 202:27 355:32]
  assign io__out_1_bits_decode_ctrl_rfWen = lsuexp | csrfix ? 1'h0 : _GEN_15; // @[SIMD_EXU.scala 357:25 358:43]
  assign io__out_1_bits_decode_ctrl_rfDest = lsuexp ? csr_bits_ctrl_rfDest : io__in_1_bits_ctrl_rfDest; // @[SIMD_EXU.scala 352:15 202:27 355:32]
  assign io__out_1_bits_decode_InstNo = lsuexp ? csr_bits_InstNo : io__in_1_bits_InstNo; // @[SIMD_EXU.scala 352:15 202:27 355:32]
  assign io__out_1_bits_decode_InstFlag = lsuexp ? csr_bits_InstFlag : io__in_1_bits_InstFlag; // @[SIMD_EXU.scala 352:15 202:27 355:32]
  assign io__out_1_bits_commits = csr_io_out_bits; // @[SIMD_EXU.scala 376:35]
  assign io__out_2_valid = SIMDU_2way_io_out_0_valid; // @[SIMD_EXU.scala 251:32]
  assign io__out_2_bits_decode_cf_pc = SIMDU_2way_io_DecodeOut_0_cf_pc; // @[SIMD_EXU.scala 247:34]
  assign io__out_2_bits_decode_cf_runahead_checkpoint_id = SIMDU_2way_io_DecodeOut_0_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 247:34]
  assign io__out_2_bits_decode_ctrl_rfWen = SIMDU_2way_io_DecodeOut_0_ctrl_rfWen; // @[SIMD_EXU.scala 249:45]
  assign io__out_2_bits_decode_ctrl_rfDest = SIMDU_2way_io_DecodeOut_0_ctrl_rfDest; // @[SIMD_EXU.scala 247:34]
  assign io__out_2_bits_decode_pext_OV = SIMDU_2way_io_DecodeOut_0_pext_OV; // @[SIMD_EXU.scala 247:34]
  assign io__out_2_bits_decode_InstNo = SIMDU_2way_io_DecodeOut_0_InstNo; // @[SIMD_EXU.scala 247:34]
  assign io__out_2_bits_commits = SIMDU_2way_io_out_0_bits; // @[SIMD_EXU.scala 253:39]
  assign io__out_3_valid = SIMDU_2way_io_out_1_valid; // @[SIMD_EXU.scala 252:33]
  assign io__out_3_bits_decode_cf_pc = SIMDU_2way_io_DecodeOut_1_cf_pc; // @[SIMD_EXU.scala 248:35]
  assign io__out_3_bits_decode_cf_runahead_checkpoint_id = SIMDU_2way_io_DecodeOut_1_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 248:35]
  assign io__out_3_bits_decode_ctrl_rfWen = SIMDU_2way_io_DecodeOut_1_ctrl_rfWen; // @[SIMD_EXU.scala 250:45]
  assign io__out_3_bits_decode_ctrl_rfDest = SIMDU_2way_io_DecodeOut_1_ctrl_rfDest; // @[SIMD_EXU.scala 248:35]
  assign io__out_3_bits_decode_pext_OV = SIMDU_2way_io_DecodeOut_1_pext_OV; // @[SIMD_EXU.scala 248:35]
  assign io__out_3_bits_decode_InstNo = SIMDU_2way_io_DecodeOut_1_InstNo; // @[SIMD_EXU.scala 248:35]
  assign io__out_3_bits_commits = SIMDU_2way_io_out_1_bits; // @[SIMD_EXU.scala 254:40]
  assign io__out_4_valid = lsu_io_out_valid & ~lsuexp; // @[SIMD_EXU.scala 370:48]
  assign io__out_4_bits_decode_cf_pc = lsu_io_DecodeOut_cf_pc; // @[SIMD_EXU.scala 309:30]
  assign io__out_4_bits_decode_cf_runahead_checkpoint_id = lsu_io_DecodeOut_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 309:30]
  assign io__out_4_bits_decode_ctrl_rfWen = lsu_io_DecodeOut_ctrl_rfWen; // @[SIMD_EXU.scala 310:41]
  assign io__out_4_bits_decode_ctrl_rfDest = lsu_io_DecodeOut_ctrl_rfDest; // @[SIMD_EXU.scala 309:30]
  assign io__out_4_bits_decode_InstNo = lsu_io_DecodeOut_InstNo; // @[SIMD_EXU.scala 309:30]
  assign io__out_4_bits_commits = lsu_io_out_bits; // @[SIMD_EXU.scala 375:35]
  assign io__out_5_valid = mdu_io_out_valid; // @[SIMD_EXU.scala 371:28]
  assign io__out_5_bits_decode_cf_pc = io__in_5_bits_cf_pc; // @[SIMD_EXU.scala 202:27]
  assign io__out_5_bits_decode_cf_runahead_checkpoint_id = io__in_5_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 202:27]
  assign io__out_5_bits_decode_ctrl_rfWen = io__in_5_bits_ctrl_rfWen; // @[SIMD_EXU.scala 203:38]
  assign io__out_5_bits_decode_ctrl_rfDest = io__in_5_bits_ctrl_rfDest; // @[SIMD_EXU.scala 202:27]
  assign io__out_5_bits_decode_InstNo = io__in_5_bits_InstNo; // @[SIMD_EXU.scala 202:27]
  assign io__out_5_bits_commits = mdu_io_out_bits; // @[SIMD_EXU.scala 377:35]
  assign io__out_6_valid = io__in_6_valid; // @[SIMD_EXU.scala 368:28]
  assign io__out_6_bits_decode_cf_pc = io__in_6_bits_cf_pc; // @[SIMD_EXU.scala 202:27]
  assign io__out_6_bits_decode_cf_redirect_target = alu_io_redirect_target; // @[SIMD_EXU.scala 365:42]
  assign io__out_6_bits_decode_cf_redirect_valid = alu_io_redirect_valid; // @[SIMD_EXU.scala 365:42]
  assign io__out_6_bits_decode_cf_runahead_checkpoint_id = io__in_6_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 202:27]
  assign io__out_6_bits_decode_ctrl_rfWen = io__in_6_bits_ctrl_rfWen; // @[SIMD_EXU.scala 203:38]
  assign io__out_6_bits_decode_ctrl_rfDest = io__in_6_bits_ctrl_rfDest; // @[SIMD_EXU.scala 202:27]
  assign io__out_6_bits_decode_InstNo = io__in_6_bits_InstNo; // @[SIMD_EXU.scala 202:27]
  assign io__out_6_bits_commits = alu_io_out_bits; // @[SIMD_EXU.scala 374:35]
  assign io__out_7_valid = io__in_7_valid; // @[SIMD_EXU.scala 369:29]
  assign io__out_7_bits_decode_cf_pc = io__in_7_bits_cf_pc; // @[SIMD_EXU.scala 202:27]
  assign io__out_7_bits_decode_cf_redirect_target = alu1_io_redirect_target; // @[SIMD_EXU.scala 366:43]
  assign io__out_7_bits_decode_cf_redirect_valid = alu1_io_redirect_valid; // @[SIMD_EXU.scala 366:43]
  assign io__out_7_bits_decode_cf_runahead_checkpoint_id = io__in_7_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 202:27]
  assign io__out_7_bits_decode_ctrl_rfWen = io__in_7_bits_ctrl_rfWen; // @[SIMD_EXU.scala 203:38]
  assign io__out_7_bits_decode_ctrl_rfDest = io__in_7_bits_ctrl_rfDest; // @[SIMD_EXU.scala 202:27]
  assign io__out_7_bits_decode_InstNo = io__in_7_bits_InstNo; // @[SIMD_EXU.scala 202:27]
  assign io__out_7_bits_commits = alu1_io_out_bits; // @[SIMD_EXU.scala 378:35]
  assign io__dmem_req_valid = lsu_io_dmem_req_valid; // @[SIMD_EXU.scala 306:11]
  assign io__dmem_req_bits_addr = lsu_io_dmem_req_bits_addr; // @[SIMD_EXU.scala 306:11]
  assign io__dmem_req_bits_size = lsu_io_dmem_req_bits_size; // @[SIMD_EXU.scala 306:11]
  assign io__dmem_req_bits_cmd = lsu_io_dmem_req_bits_cmd; // @[SIMD_EXU.scala 306:11]
  assign io__dmem_req_bits_wmask = lsu_io_dmem_req_bits_wmask; // @[SIMD_EXU.scala 306:11]
  assign io__dmem_req_bits_wdata = lsu_io_dmem_req_bits_wdata; // @[SIMD_EXU.scala 306:11]
  assign io__forward_0_valid = io__out_0_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_0_wb_rfWen = io__out_0_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_0_wb_rfDest = io__out_0_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_0_wb_rfData = io__out_0_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_0_InstNo = io__out_0_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_1_valid = io__out_1_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_1_wb_rfWen = io__out_1_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_1_wb_rfDest = io__out_1_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_1_wb_rfData = io__out_1_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_1_InstNo = io__out_1_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_2_valid = io__out_2_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_2_wb_rfWen = io__out_2_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_2_wb_rfDest = io__out_2_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_2_wb_rfData = io__out_2_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_2_InstNo = io__out_2_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_3_valid = io__out_3_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_3_wb_rfWen = io__out_3_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_3_wb_rfDest = io__out_3_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_3_wb_rfData = io__out_3_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_3_InstNo = io__out_3_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_4_valid = io__out_4_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_4_wb_rfWen = io__out_4_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_4_wb_rfDest = io__out_4_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_4_wb_rfData = io__out_4_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_4_InstNo = io__out_4_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_5_valid = io__out_5_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_5_wb_rfWen = io__out_5_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_5_wb_rfDest = io__out_5_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_5_wb_rfData = io__out_5_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_5_InstNo = io__out_5_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_6_valid = io__out_6_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_6_wb_rfWen = io__out_6_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_6_wb_rfDest = io__out_6_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_6_wb_rfData = io__out_6_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_6_InstNo = io__out_6_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__forward_7_valid = io__out_7_valid; // @[SIMD_EXU.scala 383:25]
  assign io__forward_7_wb_rfWen = io__out_7_bits_decode_ctrl_rfWen; // @[SIMD_EXU.scala 384:28]
  assign io__forward_7_wb_rfDest = io__out_7_bits_decode_ctrl_rfDest; // @[SIMD_EXU.scala 385:29]
  assign io__forward_7_wb_rfData = io__out_7_bits_commits; // @[SIMD_EXU.scala 386:29]
  assign io__forward_7_InstNo = io__out_7_bits_decode_InstNo; // @[SIMD_EXU.scala 388:26]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[SIMD_EXU.scala 349:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[SIMD_EXU.scala 350:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[SIMD_EXU.scala 350:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[SIMD_EXU.scala 350:18]
  assign lsu_firststage_fire = lsu_lsu_firststage_fire_0;
  assign flushICache = csr_flushICache_0;
  assign perfCnts_2 = PerfU_perfCnts_2_0;
  assign _WIRE_2_0 = _WIRE_2;
  assign satp = csr_satp_0;
  assign bpuUpdateReq_valid = ALU_bpuUpdateReq_0_valid;
  assign bpuUpdateReq_pc = ALU_bpuUpdateReq_0_pc;
  assign bpuUpdateReq_isMissPredict = ALU_bpuUpdateReq_0_isMissPredict;
  assign bpuUpdateReq_actualTarget = ALU_bpuUpdateReq_0_actualTarget;
  assign bpuUpdateReq_actualTaken = ALU_bpuUpdateReq_0_actualTaken;
  assign bpuUpdateReq_fuOpType = ALU_bpuUpdateReq_0_fuOpType;
  assign bpuUpdateReq_btbType = ALU_bpuUpdateReq_0_btbType;
  assign bpuUpdateReq_isRVC = ALU_bpuUpdateReq_0_isRVC;
  assign amoReq = lsu_amoReq;
  assign intrVec = csr_intrVec_0;
  assign _WIRE_1_0 = _WIRE_1;
  assign flushTLB = csr_flushTLB_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = io__in_6_valid; // @[ALU.scala 87:16]
  assign alu_io_in_bits_src1 = io__in_6_bits_data_src1; // @[SIMD_EXU.scala 190:{25,25}]
  assign alu_io_in_bits_src2 = io__in_6_bits_data_src2; // @[SIMD_EXU.scala 191:{25,25}]
  assign alu_io_in_bits_func = io__in_6_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 193:{25,25}]
  assign alu_io_cfIn_instr = io__in_6_bits_cf_instr; // @[SIMD_EXU.scala 214:15]
  assign alu_io_cfIn_pc = io__in_6_bits_cf_pc; // @[SIMD_EXU.scala 214:15]
  assign alu_io_cfIn_pnpc = io__in_6_bits_cf_pnpc; // @[SIMD_EXU.scala 214:15]
  assign alu_io_cfIn_brIdx = io__in_6_bits_cf_brIdx; // @[SIMD_EXU.scala 214:15]
  assign alu_io_offset = io__in_6_bits_data_imm; // @[SIMD_EXU.scala 215:17]
  assign alu1_clock = clock;
  assign alu1_reset = reset;
  assign alu1_io_in_valid = io__in_7_valid; // @[ALU.scala 87:16]
  assign alu1_io_in_bits_src1 = io__in_7_bits_data_src1; // @[SIMD_EXU.scala 190:{25,25}]
  assign alu1_io_in_bits_src2 = io__in_7_bits_data_src2; // @[SIMD_EXU.scala 191:{25,25}]
  assign alu1_io_in_bits_func = io__in_7_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 193:{25,25}]
  assign alu1_io_cfIn_instr = io__in_7_bits_cf_instr; // @[SIMD_EXU.scala 224:16]
  assign alu1_io_cfIn_pc = io__in_7_bits_cf_pc; // @[SIMD_EXU.scala 224:16]
  assign alu1_io_cfIn_pnpc = io__in_7_bits_cf_pnpc; // @[SIMD_EXU.scala 224:16]
  assign alu1_io_cfIn_brIdx = io__in_7_bits_cf_brIdx; // @[SIMD_EXU.scala 224:16]
  assign alu1_io_offset = io__in_7_bits_data_imm; // @[SIMD_EXU.scala 225:18]
  assign SIMDU_2way_clock = clock;
  assign SIMDU_2way_reset = reset;
  assign SIMDU_2way_io_flush = io__flush; // @[SIMD_EXU.scala 239:20]
  assign SIMDU_2way_io_DecodeIn_0_cf_instr = io__in_2_bits_cf_instr; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_cf_pc = io__in_2_bits_cf_pc; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_cf_runahead_checkpoint_id = io__in_2_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_cf_instrType = io__in_2_bits_cf_instrType; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_ctrl_fuOpType = io__in_2_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_ctrl_funct3 = io__in_2_bits_ctrl_funct3; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_ctrl_func24 = io__in_2_bits_ctrl_func24; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_ctrl_func23 = io__in_2_bits_ctrl_func23; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_ctrl_rfWen = io__in_2_bits_ctrl_rfWen; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_ctrl_rfDest = io__in_2_bits_ctrl_rfDest; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_data_src1 = io__in_2_bits_data_src1; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_data_src2 = io__in_2_bits_data_src2; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_data_src3 = io__in_2_bits_data_src3; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_InstNo = io__in_2_bits_InstNo; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_0_InstFlag = io__in_2_bits_InstFlag; // @[SIMD_EXU.scala 235:26]
  assign SIMDU_2way_io_DecodeIn_1_cf_instr = io__in_3_bits_cf_instr; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_cf_pc = io__in_3_bits_cf_pc; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_cf_runahead_checkpoint_id = io__in_3_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_cf_instrType = io__in_3_bits_cf_instrType; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_ctrl_fuOpType = io__in_3_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_ctrl_funct3 = io__in_3_bits_ctrl_funct3; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_ctrl_func24 = io__in_3_bits_ctrl_func24; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_ctrl_func23 = io__in_3_bits_ctrl_func23; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_ctrl_rfWen = io__in_3_bits_ctrl_rfWen; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_ctrl_rfDest = io__in_3_bits_ctrl_rfDest; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_data_src1 = io__in_3_bits_data_src1; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_data_src2 = io__in_3_bits_data_src2; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_data_src3 = io__in_3_bits_data_src3; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_InstNo = io__in_3_bits_InstNo; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_DecodeIn_1_InstFlag = io__in_3_bits_InstFlag; // @[SIMD_EXU.scala 236:26]
  assign SIMDU_2way_io_in_0_valid = io__in_2_valid; // @[SIMDU.scala 440:16]
  assign SIMDU_2way_io_in_1_valid = io__in_3_valid; // @[SIMDU.scala 444:16]
  assign SIMDU_2way_io_out_0_ready = io__out_2_ready; // @[SIMD_EXU.scala 237:27]
  assign SIMDU_2way_io_out_1_ready = io__out_3_ready; // @[SIMD_EXU.scala 238:27]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = io__in_5_valid; // @[MDU.scala 168:16]
  assign mdu_io_in_bits_src1 = io__in_5_bits_data_src1; // @[SIMD_EXU.scala 190:{25,25}]
  assign mdu_io_in_bits_src2 = io__in_5_bits_data_src2; // @[SIMD_EXU.scala 191:{25,25}]
  assign mdu_io_in_bits_func = io__in_5_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 193:{25,25}]
  assign mdu_io_out_ready = io__out_5_ready; // @[SIMD_EXU.scala 279:20]
  assign mdu_io_flush = io__flush; // @[SIMD_EXU.scala 280:16]
  assign ALU_clock = clock;
  assign ALU_reset = reset;
  assign ALU_io_in_valid = io__in_0_valid; // @[ALU.scala 87:16]
  assign ALU_io_in_bits_src1 = io__in_0_bits_data_src1; // @[SIMD_EXU.scala 190:{25,25}]
  assign ALU_io_in_bits_src2 = io__in_0_bits_data_src2; // @[SIMD_EXU.scala 191:{25,25}]
  assign ALU_io_in_bits_func = io__in_0_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 193:{25,25}]
  assign ALU_io_out_ready = io__out_0_ready; // @[SIMD_EXU.scala 289:22]
  assign ALU_io_cfIn_instr = io__in_0_bits_cf_instr; // @[SIMD_EXU.scala 287:17]
  assign ALU_io_cfIn_pc = io__in_0_bits_cf_pc; // @[SIMD_EXU.scala 287:17]
  assign ALU_io_cfIn_pnpc = io__in_0_bits_cf_pnpc; // @[SIMD_EXU.scala 287:17]
  assign ALU_io_cfIn_brIdx = io__in_0_bits_cf_brIdx; // @[SIMD_EXU.scala 287:17]
  assign ALU_io_offset = io__in_0_bits_data_imm; // @[SIMD_EXU.scala 288:19]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_in_valid = io__in_4_valid & ~BeforeLSUhasRedirect; // @[SIMD_EXU.scala 300:55]
  assign lsu_io_in_bits_src1 = io__in_4_bits_data_src1; // @[SIMD_EXU.scala 190:{25,25}]
  assign lsu_io_in_bits_src2 = io__in_4_bits_data_imm; // @[SIMD_PipeLSU.scala 648:15]
  assign lsu_io_in_bits_func = io__in_4_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 193:{25,25}]
  assign lsu_io_out_ready = io__out_4_ready; // @[SIMD_EXU.scala 307:20]
  assign lsu_io_wdata = io__in_4_bits_data_src2; // @[SIMD_EXU.scala 191:{25,25}]
  assign lsu_io_dmem_req_ready = io__dmem_req_ready; // @[SIMD_EXU.scala 306:11]
  assign lsu_io_dmem_resp_valid = io__dmem_resp_valid; // @[SIMD_EXU.scala 306:11]
  assign lsu_io_dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[SIMD_EXU.scala 306:11]
  assign lsu_io_flush = io__flush; // @[SIMD_EXU.scala 308:16]
  assign lsu_io_DecodeIn_cf_instr = io__in_4_bits_cf_instr; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_pc = io__in_4_bits_cf_pc; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_exceptionVec_1 = io__in_4_bits_cf_exceptionVec_1; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_exceptionVec_2 = io__in_4_bits_cf_exceptionVec_2; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_exceptionVec_12 = io__in_4_bits_cf_exceptionVec_12; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_0 = io__in_4_bits_cf_intrVec_0; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_1 = io__in_4_bits_cf_intrVec_1; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_2 = io__in_4_bits_cf_intrVec_2; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_3 = io__in_4_bits_cf_intrVec_3; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_4 = io__in_4_bits_cf_intrVec_4; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_5 = io__in_4_bits_cf_intrVec_5; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_6 = io__in_4_bits_cf_intrVec_6; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_7 = io__in_4_bits_cf_intrVec_7; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_8 = io__in_4_bits_cf_intrVec_8; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_9 = io__in_4_bits_cf_intrVec_9; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_10 = io__in_4_bits_cf_intrVec_10; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_intrVec_11 = io__in_4_bits_cf_intrVec_11; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_crossPageIPFFix = io__in_4_bits_cf_crossPageIPFFix; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_cf_runahead_checkpoint_id = io__in_4_bits_cf_runahead_checkpoint_id; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_ctrl_rfWen = io__in_4_bits_ctrl_rfWen; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_ctrl_rfDest = io__in_4_bits_ctrl_rfDest; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_ctrl_isMou = io__in_4_bits_ctrl_isMou; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_InstNo = io__in_4_bits_InstNo; // @[SIMD_EXU.scala 299:19]
  assign lsu_io_DecodeIn_InstFlag = io__in_4_bits_InstFlag; // @[SIMD_EXU.scala 299:19]
  assign lsu__T_408 = _T_408;
  assign lsu_io_memMMU_dmem_loadPF = io__memMMU_dmem_loadPF;
  assign lsu_ismmio = ismmio;
  assign lsu_lr = csr_lr_0;
  assign lsu_io_memMMU_dmem_storePF = io__memMMU_dmem_storePF;
  assign lsu_vmEnable = vmEnable;
  assign lsu__T_407 = _T_407;
  assign lsu_lrAddr = csr_lrAddr_0;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = io__in_1_valid; // @[SIMD_CSR.scala 504:16]
  assign csr_io_in_bits_src1 = io__in_1_bits_data_src1; // @[SIMD_EXU.scala 190:{25,25}]
  assign csr_io_in_bits_src2 = io__in_1_bits_data_src2; // @[SIMD_EXU.scala 191:{25,25}]
  assign csr_io_in_bits_func = io__in_1_bits_ctrl_fuOpType; // @[SIMD_EXU.scala 193:{25,25}]
  assign csr_io_cfIn_pc = io__in_1_valid ? io__in_1_bits_cf_pc : lsu_io_DecodeOut_cf_pc; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_exceptionVec_1 = io__in_1_valid ? io__in_1_bits_cf_exceptionVec_1 :
    lsu_io_DecodeOut_cf_exceptionVec_1; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_exceptionVec_2 = io__in_1_valid ? io__in_1_bits_cf_exceptionVec_2 :
    lsu_io_DecodeOut_cf_exceptionVec_2; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io_loadAddrMisaligned; // @[SIMD_EXU.scala 320:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io_storeAddrMisaligned; // @[SIMD_EXU.scala 321:49]
  assign csr_io_cfIn_exceptionVec_12 = io__in_1_valid ? io__in_1_bits_cf_exceptionVec_12 :
    lsu_io_DecodeOut_cf_exceptionVec_12; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_exceptionVec_13 = lsu_io_loadPF; // @[SIMD_EXU.scala 338:43]
  assign csr_io_cfIn_exceptionVec_15 = lsu_io_storePF; // @[SIMD_EXU.scala 339:44]
  assign csr_io_cfIn_intrVec_0 = io__in_1_valid ? io__in_1_bits_cf_intrVec_0 : lsu_io_DecodeOut_cf_intrVec_0; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_1 = io__in_1_valid ? io__in_1_bits_cf_intrVec_1 : lsu_io_DecodeOut_cf_intrVec_1; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_2 = io__in_1_valid ? io__in_1_bits_cf_intrVec_2 : lsu_io_DecodeOut_cf_intrVec_2; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_3 = io__in_1_valid ? io__in_1_bits_cf_intrVec_3 : lsu_io_DecodeOut_cf_intrVec_3; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_4 = io__in_1_valid ? io__in_1_bits_cf_intrVec_4 : lsu_io_DecodeOut_cf_intrVec_4; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_5 = io__in_1_valid ? io__in_1_bits_cf_intrVec_5 : lsu_io_DecodeOut_cf_intrVec_5; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_6 = io__in_1_valid ? io__in_1_bits_cf_intrVec_6 : lsu_io_DecodeOut_cf_intrVec_6; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_7 = io__in_1_valid ? io__in_1_bits_cf_intrVec_7 : lsu_io_DecodeOut_cf_intrVec_7; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_8 = io__in_1_valid ? io__in_1_bits_cf_intrVec_8 : lsu_io_DecodeOut_cf_intrVec_8; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_9 = io__in_1_valid ? io__in_1_bits_cf_intrVec_9 : lsu_io_DecodeOut_cf_intrVec_9; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_10 = io__in_1_valid ? io__in_1_bits_cf_intrVec_10 : lsu_io_DecodeOut_cf_intrVec_10; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_intrVec_11 = io__in_1_valid ? io__in_1_bits_cf_intrVec_11 : lsu_io_DecodeOut_cf_intrVec_11; // @[SIMD_EXU.scala 318:21]
  assign csr_io_cfIn_crossPageIPFFix = io__in_1_valid ? io__in_1_bits_cf_crossPageIPFFix :
    lsu_io_DecodeOut_cf_crossPageIPFFix; // @[SIMD_EXU.scala 318:21]
  assign csr_io_ctrlIn_isMou = io__in_1_valid ? io__in_1_bits_ctrl_isMou : lsu_io_DecodeOut_ctrl_isMou; // @[SIMD_EXU.scala 319:23]
  assign csr_io_instrValid = (io__in_1_valid | lsuexp) & _T_4; // @[SIMD_EXU.scala 342:56]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[SIMD_EXU.scala 350:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[SIMD_EXU.scala 350:18]
  assign csr_io_dmemMMU_addr = io__memMMU_dmem_addr; // @[SIMD_EXU.scala 350:18]
  assign csr_set_lr = lsu_setLr;
  assign csr_OVWEN_0 = _WIRE_2_1;
  assign csr_mtip = io_extra_mtip;
  assign csr_meip = io_extra_meip_0;
  assign csr_LSUADDR = lsu_addr_0;
  assign csr_msip = io_extra_msip;
  assign csr_set_lr_addr = lsu_setLrAddr;
  assign csr_set_lr_val = lsu_setLrVal;
  assign PerfU_clock = clock;
  assign PerfU_reset = reset;
  assign PerfU_perfCntCondMultiCommit3 = _T_137_0;
  assign PerfU_perfCntCondMultiCommit6 = _T_140_0;
  assign PerfU_perfCntCondMinstret = io_in_0_valid;
  assign PerfU_perfCntCondMultiCommit2 = _T_136_0;
  assign PerfU_perfCntCondMultiCommit5 = _T_139_0;
  assign PerfU_perfCntCondMultiCommit4 = _T_138_0;
  assign PerfU_perfCntCondMultiCommit = _T_135_0;
endmodule
module new_SIMD_WBU(
  input         clock,
  input         reset,
  input         io__in_0_valid,
  input  [38:0] io__in_0_bits_decode_cf_pc,
  input  [38:0] io__in_0_bits_decode_cf_redirect_target,
  input         io__in_0_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_0_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_0_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_0_bits_decode_ctrl_rfDest,
  input         io__in_0_bits_decode_pext_OV,
  input  [4:0]  io__in_0_bits_decode_InstNo,
  input  [63:0] io__in_0_bits_commits,
  input         io__in_1_valid,
  input  [38:0] io__in_1_bits_decode_cf_pc,
  input  [38:0] io__in_1_bits_decode_cf_redirect_target,
  input         io__in_1_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_1_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_1_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_1_bits_decode_ctrl_rfDest,
  input         io__in_1_bits_decode_pext_OV,
  input  [4:0]  io__in_1_bits_decode_InstNo,
  input  [63:0] io__in_1_bits_commits,
  input         io__in_2_valid,
  input  [38:0] io__in_2_bits_decode_cf_pc,
  input  [38:0] io__in_2_bits_decode_cf_redirect_target,
  input         io__in_2_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_2_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_2_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_2_bits_decode_ctrl_rfDest,
  input         io__in_2_bits_decode_pext_OV,
  input  [4:0]  io__in_2_bits_decode_InstNo,
  input  [63:0] io__in_2_bits_commits,
  input         io__in_3_valid,
  input  [38:0] io__in_3_bits_decode_cf_pc,
  input  [38:0] io__in_3_bits_decode_cf_redirect_target,
  input         io__in_3_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_3_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_3_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_3_bits_decode_ctrl_rfDest,
  input         io__in_3_bits_decode_pext_OV,
  input  [4:0]  io__in_3_bits_decode_InstNo,
  input  [63:0] io__in_3_bits_commits,
  input         io__in_4_valid,
  input  [38:0] io__in_4_bits_decode_cf_pc,
  input  [38:0] io__in_4_bits_decode_cf_redirect_target,
  input         io__in_4_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_4_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_4_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_4_bits_decode_ctrl_rfDest,
  input         io__in_4_bits_decode_pext_OV,
  input  [4:0]  io__in_4_bits_decode_InstNo,
  input  [63:0] io__in_4_bits_commits,
  input         io__in_5_valid,
  input  [38:0] io__in_5_bits_decode_cf_pc,
  input  [38:0] io__in_5_bits_decode_cf_redirect_target,
  input         io__in_5_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_5_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_5_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_5_bits_decode_ctrl_rfDest,
  input         io__in_5_bits_decode_pext_OV,
  input  [4:0]  io__in_5_bits_decode_InstNo,
  input  [63:0] io__in_5_bits_commits,
  input         io__in_6_valid,
  input  [38:0] io__in_6_bits_decode_cf_pc,
  input  [38:0] io__in_6_bits_decode_cf_redirect_target,
  input         io__in_6_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_6_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_6_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_6_bits_decode_ctrl_rfDest,
  input         io__in_6_bits_decode_pext_OV,
  input  [4:0]  io__in_6_bits_decode_InstNo,
  input  [63:0] io__in_6_bits_commits,
  input         io__in_7_valid,
  input  [38:0] io__in_7_bits_decode_cf_pc,
  input  [38:0] io__in_7_bits_decode_cf_redirect_target,
  input         io__in_7_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_7_bits_decode_cf_runahead_checkpoint_id,
  input         io__in_7_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_7_bits_decode_ctrl_rfDest,
  input         io__in_7_bits_decode_pext_OV,
  input  [4:0]  io__in_7_bits_decode_InstNo,
  input  [63:0] io__in_7_bits_commits,
  output        io__wb_rfWen_0,
  output        io__wb_rfWen_1,
  output        io__wb_rfWen_2,
  output        io__wb_rfWen_3,
  output        io__wb_rfWen_4,
  output        io__wb_rfWen_5,
  output        io__wb_rfWen_6,
  output        io__wb_rfWen_7,
  output [4:0]  io__wb_rfDest_0,
  output [4:0]  io__wb_rfDest_1,
  output [4:0]  io__wb_rfDest_2,
  output [4:0]  io__wb_rfDest_3,
  output [4:0]  io__wb_rfDest_4,
  output [4:0]  io__wb_rfDest_5,
  output [4:0]  io__wb_rfDest_6,
  output [4:0]  io__wb_rfDest_7,
  output [63:0] io__wb_WriteData_0,
  output [63:0] io__wb_WriteData_1,
  output [63:0] io__wb_WriteData_2,
  output [63:0] io__wb_WriteData_3,
  output [63:0] io__wb_WriteData_4,
  output [63:0] io__wb_WriteData_5,
  output [63:0] io__wb_WriteData_6,
  output [63:0] io__wb_WriteData_7,
  input  [4:0]  io__wb_rfSrc1_0,
  input  [4:0]  io__wb_rfSrc1_1,
  input  [4:0]  io__wb_rfSrc2_0,
  input  [4:0]  io__wb_rfSrc2_1,
  input  [4:0]  io__wb_rfSrc3_0,
  input  [4:0]  io__wb_rfSrc3_1,
  output [63:0] io__wb_ReadData1_0,
  output [63:0] io__wb_ReadData1_1,
  output [63:0] io__wb_ReadData2_0,
  output [63:0] io__wb_ReadData2_1,
  output [63:0] io__wb_ReadData3_0,
  output [63:0] io__wb_ReadData3_1,
  output [4:0]  io__wb_InstNo_0,
  output [4:0]  io__wb_InstNo_1,
  output [4:0]  io__wb_InstNo_2,
  output [4:0]  io__wb_InstNo_3,
  output [4:0]  io__wb_InstNo_4,
  output [4:0]  io__wb_InstNo_5,
  output [4:0]  io__wb_InstNo_6,
  output [4:0]  io__wb_InstNo_7,
  output        io__redirect_valid,
  output        _T_137_0,
  output        _T_140_0,
  output [38:0] io_in_0_bits_decode_cf_pc,
  output [4:0]  io_wb_rfDest_0,
  output        io_in_0_valid,
  output        _WIRE_2_1,
  output        _T_136_0,
  output        _T_139_0,
  output        io_wb_rfWen_0,
  output [63:0] io_wb_WriteData_0,
  output        _T_138_0,
  output        io_in_0_valid_0,
  output        _T_135_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] MEM [0:31]; // @[RF.scala 31:15]
  wire  MEM_MPORT_16_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_16_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_16_data; // @[RF.scala 31:15]
  wire  MEM_MPORT_17_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_17_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_17_data; // @[RF.scala 31:15]
  wire  MEM_MPORT_18_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_18_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_18_data; // @[RF.scala 31:15]
  wire  MEM_MPORT_19_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_19_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_19_data; // @[RF.scala 31:15]
  wire  MEM_MPORT_20_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_20_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_20_data; // @[RF.scala 31:15]
  wire  MEM_MPORT_21_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_21_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_21_data; // @[RF.scala 31:15]
  wire  MEM_MPORT_22_en; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_22_addr; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_22_data; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_1_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_1_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_1_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_1_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_2_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_2_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_2_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_2_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_3_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_3_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_3_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_3_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_4_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_4_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_4_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_4_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_5_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_5_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_5_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_5_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_6_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_6_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_6_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_6_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_7_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_7_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_7_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_7_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_8_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_8_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_8_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_8_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_9_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_9_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_9_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_9_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_10_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_10_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_10_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_10_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_11_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_11_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_11_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_11_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_12_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_12_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_12_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_12_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_13_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_13_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_13_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_13_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_14_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_14_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_14_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_14_en; // @[RF.scala 31:15]
  wire [63:0] MEM_MPORT_15_data; // @[RF.scala 31:15]
  wire [4:0] MEM_MPORT_15_addr; // @[RF.scala 31:15]
  wire  MEM_MPORT_15_mask; // @[RF.scala 31:15]
  wire  MEM_MPORT_15_en; // @[RF.scala 31:15]
  wire  runahead_redirect_io_clock; // @[SIMD_WBU.scala 167:33]
  wire [7:0] runahead_redirect_io_coreid; // @[SIMD_WBU.scala 167:33]
  wire  runahead_redirect_io_valid; // @[SIMD_WBU.scala 167:33]
  wire [63:0] runahead_redirect_io_pc; // @[SIMD_WBU.scala 167:33]
  wire [63:0] runahead_redirect_io_target_pc; // @[SIMD_WBU.scala 167:33]
  wire [63:0] runahead_redirect_io_checkpoint_id; // @[SIMD_WBU.scala 167:33]
  wire  _T = io__in_0_bits_decode_cf_redirect_valid & io__in_0_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_1 = io__in_1_bits_decode_cf_redirect_valid & io__in_1_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_2 = io__in_2_bits_decode_cf_redirect_valid & io__in_2_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_3 = io__in_3_bits_decode_cf_redirect_valid & io__in_3_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_4 = io__in_4_bits_decode_cf_redirect_valid & io__in_4_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_5 = io__in_5_bits_decode_cf_redirect_valid & io__in_5_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_6 = io__in_6_bits_decode_cf_redirect_valid & io__in_6_valid; // @[SIMD_WBU.scala 127:111]
  wire  _T_7 = io__in_7_bits_decode_cf_redirect_valid & io__in_7_valid; // @[SIMD_WBU.scala 127:111]
  wire [2:0] _T_8 = _T_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_9 = _T_5 ? 3'h5 : _T_8; // @[Mux.scala 47:69]
  wire [2:0] _T_10 = _T_4 ? 3'h4 : _T_9; // @[Mux.scala 47:69]
  wire [2:0] _T_11 = _T_3 ? 3'h3 : _T_10; // @[Mux.scala 47:69]
  wire [2:0] _T_12 = _T_2 ? 3'h2 : _T_11; // @[Mux.scala 47:69]
  wire [2:0] _T_13 = _T_1 ? 3'h1 : _T_12; // @[Mux.scala 47:69]
  wire [2:0] redirct_index = _T ? 3'h0 : _T_13; // @[Mux.scala 47:69]
  wire [38:0] _GEN_17 = 3'h1 == redirct_index ? io__in_1_bits_decode_cf_redirect_target :
    io__in_0_bits_decode_cf_redirect_target; // @[SIMD_WBU.scala 128:{15,15}]
  wire [38:0] _GEN_18 = 3'h2 == redirct_index ? io__in_2_bits_decode_cf_redirect_target : _GEN_17; // @[SIMD_WBU.scala 128:{15,15}]
  wire [38:0] _GEN_19 = 3'h3 == redirct_index ? io__in_3_bits_decode_cf_redirect_target : _GEN_18; // @[SIMD_WBU.scala 128:{15,15}]
  wire [38:0] _GEN_20 = 3'h4 == redirct_index ? io__in_4_bits_decode_cf_redirect_target : _GEN_19; // @[SIMD_WBU.scala 128:{15,15}]
  wire [38:0] _GEN_21 = 3'h5 == redirct_index ? io__in_5_bits_decode_cf_redirect_target : _GEN_20; // @[SIMD_WBU.scala 128:{15,15}]
  wire [38:0] _GEN_22 = 3'h6 == redirct_index ? io__in_6_bits_decode_cf_redirect_target : _GEN_21; // @[SIMD_WBU.scala 128:{15,15}]
  wire [38:0] _GEN_23 = 3'h7 == redirct_index ? io__in_7_bits_decode_cf_redirect_target : _GEN_22; // @[SIMD_WBU.scala 128:{15,15}]
  wire  FronthasRedirect_1 = 3'h1 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  FronthasRedirect_2 = 3'h2 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  FronthasRedirect_3 = 3'h3 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  FronthasRedirect_4 = 3'h4 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  FronthasRedirect_5 = 3'h5 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  FronthasRedirect_6 = 3'h6 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  FronthasRedirect_7 = 3'h7 > redirct_index; // @[SIMD_WBU.scala 131:67]
  wire  _T_49 = ~FronthasRedirect_1; // @[SIMD_WBU.scala 141:29]
  wire  _T_53 = ~FronthasRedirect_2; // @[SIMD_WBU.scala 141:29]
  wire  _T_57 = ~FronthasRedirect_3; // @[SIMD_WBU.scala 141:29]
  wire  _T_61 = ~FronthasRedirect_4; // @[SIMD_WBU.scala 141:29]
  wire  _T_65 = ~FronthasRedirect_5; // @[SIMD_WBU.scala 141:29]
  wire  _T_69 = ~FronthasRedirect_6; // @[SIMD_WBU.scala 141:29]
  wire  _T_73 = ~FronthasRedirect_7; // @[SIMD_WBU.scala 141:29]
  wire [38:0] _GEN_113 = 3'h1 == redirct_index ? io__in_1_bits_decode_cf_pc : io__in_0_bits_decode_cf_pc; // @[SIMD_WBU.scala 171:{27,27}]
  wire [38:0] _GEN_114 = 3'h2 == redirct_index ? io__in_2_bits_decode_cf_pc : _GEN_113; // @[SIMD_WBU.scala 171:{27,27}]
  wire [38:0] _GEN_115 = 3'h3 == redirct_index ? io__in_3_bits_decode_cf_pc : _GEN_114; // @[SIMD_WBU.scala 171:{27,27}]
  wire [38:0] _GEN_116 = 3'h4 == redirct_index ? io__in_4_bits_decode_cf_pc : _GEN_115; // @[SIMD_WBU.scala 171:{27,27}]
  wire [38:0] _GEN_117 = 3'h5 == redirct_index ? io__in_5_bits_decode_cf_pc : _GEN_116; // @[SIMD_WBU.scala 171:{27,27}]
  wire [38:0] _GEN_118 = 3'h6 == redirct_index ? io__in_6_bits_decode_cf_pc : _GEN_117; // @[SIMD_WBU.scala 171:{27,27}]
  wire [38:0] _GEN_119 = 3'h7 == redirct_index ? io__in_7_bits_decode_cf_pc : _GEN_118; // @[SIMD_WBU.scala 171:{27,27}]
  wire [63:0] _GEN_121 = 3'h1 == redirct_index ? io__in_1_bits_decode_cf_runahead_checkpoint_id :
    io__in_0_bits_decode_cf_runahead_checkpoint_id; // @[SIMD_WBU.scala 173:{38,38}]
  wire [63:0] _GEN_122 = 3'h2 == redirct_index ? io__in_2_bits_decode_cf_runahead_checkpoint_id : _GEN_121; // @[SIMD_WBU.scala 173:{38,38}]
  wire [63:0] _GEN_123 = 3'h3 == redirct_index ? io__in_3_bits_decode_cf_runahead_checkpoint_id : _GEN_122; // @[SIMD_WBU.scala 173:{38,38}]
  wire [63:0] _GEN_124 = 3'h4 == redirct_index ? io__in_4_bits_decode_cf_runahead_checkpoint_id : _GEN_123; // @[SIMD_WBU.scala 173:{38,38}]
  wire [63:0] _GEN_125 = 3'h5 == redirct_index ? io__in_5_bits_decode_cf_runahead_checkpoint_id : _GEN_124; // @[SIMD_WBU.scala 173:{38,38}]
  wire [63:0] _GEN_126 = 3'h6 == redirct_index ? io__in_6_bits_decode_cf_runahead_checkpoint_id : _GEN_125; // @[SIMD_WBU.scala 173:{38,38}]
  wire  _T_116 = io__in_1_valid & _T_49; // @[SIMD_WBU.scala 178:65]
  wire  _T_118 = io__in_2_valid & _T_53; // @[SIMD_WBU.scala 178:65]
  wire  _T_120 = io__in_3_valid & _T_57; // @[SIMD_WBU.scala 178:65]
  wire  _T_122 = io__in_4_valid & _T_61; // @[SIMD_WBU.scala 178:65]
  wire  _T_124 = io__in_5_valid & _T_65; // @[SIMD_WBU.scala 178:65]
  wire  _T_126 = io__in_6_valid & _T_69; // @[SIMD_WBU.scala 178:65]
  wire  _T_128 = io__in_7_valid & _T_73; // @[SIMD_WBU.scala 178:65]
  wire [1:0] _T_129 = io__in_0_valid + _T_116; // @[SIMD_WBU.scala 178:106]
  wire [1:0] _GEN_128 = {{1'd0}, _T_118}; // @[SIMD_WBU.scala 178:106]
  wire [2:0] _T_130 = _T_129 + _GEN_128; // @[SIMD_WBU.scala 178:106]
  wire [2:0] _GEN_129 = {{2'd0}, _T_120}; // @[SIMD_WBU.scala 178:106]
  wire [3:0] _T_131 = _T_130 + _GEN_129; // @[SIMD_WBU.scala 178:106]
  wire [3:0] _GEN_130 = {{3'd0}, _T_122}; // @[SIMD_WBU.scala 178:106]
  wire [4:0] _T_132 = _T_131 + _GEN_130; // @[SIMD_WBU.scala 178:106]
  wire [4:0] _GEN_131 = {{4'd0}, _T_124}; // @[SIMD_WBU.scala 178:106]
  wire [5:0] _T_133 = _T_132 + _GEN_131; // @[SIMD_WBU.scala 178:106]
  wire [5:0] _GEN_132 = {{5'd0}, _T_126}; // @[SIMD_WBU.scala 178:106]
  wire [6:0] _T_134 = _T_133 + _GEN_132; // @[SIMD_WBU.scala 178:106]
  wire [6:0] _GEN_133 = {{6'd0}, _T_128}; // @[SIMD_WBU.scala 178:106]
  wire [7:0] commit_num = _T_134 + _GEN_133; // @[SIMD_WBU.scala 178:106]
  wire  _T_135 = commit_num != 8'h0; // @[SIMD_WBU.scala 181:35]
  wire  _T_136 = commit_num == 8'h2; // @[SIMD_WBU.scala 182:35]
  wire  _T_137 = commit_num == 8'h3; // @[SIMD_WBU.scala 183:35]
  wire  _T_138 = commit_num == 8'h4; // @[SIMD_WBU.scala 184:35]
  wire  _T_139 = commit_num == 8'h5; // @[SIMD_WBU.scala 185:35]
  wire  _T_140 = commit_num == 8'h6; // @[SIMD_WBU.scala 186:35]
  wire  _WIRE_2 = io__in_7_valid & io__in_7_bits_decode_pext_OV & _T_73 | (io__in_6_valid & io__in_6_bits_decode_pext_OV
     & _T_69 | (io__in_5_valid & io__in_5_bits_decode_pext_OV & _T_65 | (io__in_4_valid & io__in_4_bits_decode_pext_OV
     & _T_61 | (io__in_3_valid & io__in_3_bits_decode_pext_OV & _T_57 | (io__in_2_valid & io__in_2_bits_decode_pext_OV
     & _T_53 | (io__in_1_valid & io__in_1_bits_decode_pext_OV & _T_49 | io__in_0_valid & io__in_0_bits_decode_pext_OV)))
    ))); // @[SIMD_WBU.scala 160:83 161:19]
  DifftestRunaheadRedirectEvent runahead_redirect ( // @[SIMD_WBU.scala 167:33]
    .io_clock(runahead_redirect_io_clock),
    .io_coreid(runahead_redirect_io_coreid),
    .io_valid(runahead_redirect_io_valid),
    .io_pc(runahead_redirect_io_pc),
    .io_target_pc(runahead_redirect_io_target_pc),
    .io_checkpoint_id(runahead_redirect_io_checkpoint_id)
  );
  assign MEM_MPORT_16_en = 1'h1;
  assign MEM_MPORT_16_addr = io__wb_rfSrc1_0;
  assign MEM_MPORT_16_data = MEM[MEM_MPORT_16_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_17_en = 1'h1;
  assign MEM_MPORT_17_addr = io__wb_rfSrc2_0;
  assign MEM_MPORT_17_data = MEM[MEM_MPORT_17_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_18_en = 1'h1;
  assign MEM_MPORT_18_addr = io__wb_rfSrc3_0;
  assign MEM_MPORT_18_data = MEM[MEM_MPORT_18_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_19_en = 1'h1;
  assign MEM_MPORT_19_addr = io__wb_rfSrc1_1;
  assign MEM_MPORT_19_data = MEM[MEM_MPORT_19_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_20_en = 1'h1;
  assign MEM_MPORT_20_addr = io__wb_rfSrc2_1;
  assign MEM_MPORT_20_data = MEM[MEM_MPORT_20_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_21_en = 1'h1;
  assign MEM_MPORT_21_addr = io__wb_rfSrc3_1;
  assign MEM_MPORT_21_data = MEM[MEM_MPORT_21_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_22_en = 1'h1;
  assign MEM_MPORT_22_addr = 5'h5;
  assign MEM_MPORT_22_data = MEM[MEM_MPORT_22_addr]; // @[RF.scala 31:15]
  assign MEM_MPORT_data = io__wb_WriteData_0;
  assign MEM_MPORT_addr = io__wb_rfDest_0;
  assign MEM_MPORT_mask = 1'h1;
  assign MEM_MPORT_en = io__wb_rfWen_0;
  assign MEM_MPORT_1_data = 64'h0;
  assign MEM_MPORT_1_addr = io__wb_rfDest_0;
  assign MEM_MPORT_1_mask = 1'h1;
  assign MEM_MPORT_1_en = reset;
  assign MEM_MPORT_2_data = io__wb_WriteData_1;
  assign MEM_MPORT_2_addr = io__wb_rfDest_1;
  assign MEM_MPORT_2_mask = 1'h1;
  assign MEM_MPORT_2_en = io__wb_rfWen_1 & _T_49;
  assign MEM_MPORT_3_data = 64'h0;
  assign MEM_MPORT_3_addr = io__wb_rfDest_1;
  assign MEM_MPORT_3_mask = 1'h1;
  assign MEM_MPORT_3_en = reset;
  assign MEM_MPORT_4_data = io__wb_WriteData_2;
  assign MEM_MPORT_4_addr = io__wb_rfDest_2;
  assign MEM_MPORT_4_mask = 1'h1;
  assign MEM_MPORT_4_en = io__wb_rfWen_2 & _T_53;
  assign MEM_MPORT_5_data = 64'h0;
  assign MEM_MPORT_5_addr = io__wb_rfDest_2;
  assign MEM_MPORT_5_mask = 1'h1;
  assign MEM_MPORT_5_en = reset;
  assign MEM_MPORT_6_data = io__wb_WriteData_3;
  assign MEM_MPORT_6_addr = io__wb_rfDest_3;
  assign MEM_MPORT_6_mask = 1'h1;
  assign MEM_MPORT_6_en = io__wb_rfWen_3 & _T_57;
  assign MEM_MPORT_7_data = 64'h0;
  assign MEM_MPORT_7_addr = io__wb_rfDest_3;
  assign MEM_MPORT_7_mask = 1'h1;
  assign MEM_MPORT_7_en = reset;
  assign MEM_MPORT_8_data = io__wb_WriteData_4;
  assign MEM_MPORT_8_addr = io__wb_rfDest_4;
  assign MEM_MPORT_8_mask = 1'h1;
  assign MEM_MPORT_8_en = io__wb_rfWen_4 & _T_61;
  assign MEM_MPORT_9_data = 64'h0;
  assign MEM_MPORT_9_addr = io__wb_rfDest_4;
  assign MEM_MPORT_9_mask = 1'h1;
  assign MEM_MPORT_9_en = reset;
  assign MEM_MPORT_10_data = io__wb_WriteData_5;
  assign MEM_MPORT_10_addr = io__wb_rfDest_5;
  assign MEM_MPORT_10_mask = 1'h1;
  assign MEM_MPORT_10_en = io__wb_rfWen_5 & _T_65;
  assign MEM_MPORT_11_data = 64'h0;
  assign MEM_MPORT_11_addr = io__wb_rfDest_5;
  assign MEM_MPORT_11_mask = 1'h1;
  assign MEM_MPORT_11_en = reset;
  assign MEM_MPORT_12_data = io__wb_WriteData_6;
  assign MEM_MPORT_12_addr = io__wb_rfDest_6;
  assign MEM_MPORT_12_mask = 1'h1;
  assign MEM_MPORT_12_en = io__wb_rfWen_6 & _T_69;
  assign MEM_MPORT_13_data = 64'h0;
  assign MEM_MPORT_13_addr = io__wb_rfDest_6;
  assign MEM_MPORT_13_mask = 1'h1;
  assign MEM_MPORT_13_en = reset;
  assign MEM_MPORT_14_data = io__wb_WriteData_7;
  assign MEM_MPORT_14_addr = io__wb_rfDest_7;
  assign MEM_MPORT_14_mask = 1'h1;
  assign MEM_MPORT_14_en = io__wb_rfWen_7 & _T_73;
  assign MEM_MPORT_15_data = 64'h0;
  assign MEM_MPORT_15_addr = io__wb_rfDest_7;
  assign MEM_MPORT_15_mask = 1'h1;
  assign MEM_MPORT_15_en = reset;
  assign io__wb_rfWen_0 = io__in_0_bits_decode_ctrl_rfWen & io__in_0_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_1 = io__in_1_bits_decode_ctrl_rfWen & io__in_1_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_2 = io__in_2_bits_decode_ctrl_rfWen & io__in_2_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_3 = io__in_3_bits_decode_ctrl_rfWen & io__in_3_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_4 = io__in_4_bits_decode_ctrl_rfWen & io__in_4_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_5 = io__in_5_bits_decode_ctrl_rfWen & io__in_5_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_6 = io__in_6_bits_decode_ctrl_rfWen & io__in_6_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfWen_7 = io__in_7_bits_decode_ctrl_rfWen & io__in_7_valid; // @[SIMD_WBU.scala 134:55]
  assign io__wb_rfDest_0 = io__in_0_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_1 = io__in_1_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_2 = io__in_2_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_3 = io__in_3_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_4 = io__in_4_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_5 = io__in_5_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_6 = io__in_6_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_rfDest_7 = io__in_7_bits_decode_ctrl_rfDest; // @[SIMD_WBU.scala 135:21]
  assign io__wb_WriteData_0 = io__in_0_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_1 = io__in_1_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_2 = io__in_2_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_3 = io__in_3_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_4 = io__in_4_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_5 = io__in_5_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_6 = io__in_6_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_WriteData_7 = io__in_7_bits_commits; // @[SIMD_WBU.scala 136:24]
  assign io__wb_ReadData1_0 = io__wb_rfSrc1_0 == 5'h0 ? 64'h0 : MEM_MPORT_16_data; // @[RF.scala 32:36]
  assign io__wb_ReadData1_1 = io__wb_rfSrc1_1 == 5'h0 ? 64'h0 : MEM_MPORT_19_data; // @[RF.scala 32:36]
  assign io__wb_ReadData2_0 = io__wb_rfSrc2_0 == 5'h0 ? 64'h0 : MEM_MPORT_17_data; // @[RF.scala 32:36]
  assign io__wb_ReadData2_1 = io__wb_rfSrc2_1 == 5'h0 ? 64'h0 : MEM_MPORT_20_data; // @[RF.scala 32:36]
  assign io__wb_ReadData3_0 = io__wb_rfSrc3_0 == 5'h0 ? 64'h0 : MEM_MPORT_18_data; // @[RF.scala 32:36]
  assign io__wb_ReadData3_1 = io__wb_rfSrc3_1 == 5'h0 ? 64'h0 : MEM_MPORT_21_data; // @[RF.scala 32:36]
  assign io__wb_InstNo_0 = io__in_0_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_1 = io__in_1_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_2 = io__in_2_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_3 = io__in_3_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_4 = io__in_4_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_5 = io__in_5_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_6 = io__in_6_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__wb_InstNo_7 = io__in_7_bits_decode_InstNo; // @[SIMD_WBU.scala 138:21]
  assign io__redirect_valid = _T | _T_1 | _T_2 | _T_3 | _T_4 | _T_5 | _T_6 | _T_7; // @[SIMD_WBU.scala 129:128]
  assign _T_137_0 = _T_137;
  assign _T_140_0 = _T_140;
  assign io_in_0_bits_decode_cf_pc = io__in_0_bits_decode_cf_pc;
  assign io_wb_rfDest_0 = io__wb_rfDest_0;
  assign io_in_0_valid = io__in_0_valid;
  assign _WIRE_2_1 = _WIRE_2;
  assign _T_136_0 = _T_136;
  assign _T_139_0 = _T_139;
  assign io_wb_rfWen_0 = io__wb_rfWen_0;
  assign io_wb_WriteData_0 = io__wb_WriteData_0;
  assign _T_138_0 = _T_138;
  assign io_in_0_valid_0 = io__in_0_valid;
  assign _T_135_0 = _T_135;
  assign runahead_redirect_io_clock = clock; // @[SIMD_WBU.scala 168:30]
  assign runahead_redirect_io_coreid = 8'h0; // @[SIMD_WBU.scala 169:31]
  assign runahead_redirect_io_valid = io__redirect_valid; // @[SIMD_WBU.scala 170:30]
  assign runahead_redirect_io_pc = {{25'd0}, _GEN_119}; // @[SIMD_WBU.scala 171:27]
  assign runahead_redirect_io_target_pc = {{25'd0}, _GEN_23}; // @[SIMD_WBU.scala 172:34]
  assign runahead_redirect_io_checkpoint_id = 3'h7 == redirct_index ? io__in_7_bits_decode_cf_runahead_checkpoint_id :
    _GEN_126; // @[SIMD_WBU.scala 173:{38,38}]
  always @(posedge clock) begin
    if (MEM_MPORT_en & MEM_MPORT_mask) begin
      MEM[MEM_MPORT_addr] <= MEM_MPORT_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_1_en & MEM_MPORT_1_mask) begin
      MEM[MEM_MPORT_1_addr] <= MEM_MPORT_1_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_2_en & MEM_MPORT_2_mask) begin
      MEM[MEM_MPORT_2_addr] <= MEM_MPORT_2_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_3_en & MEM_MPORT_3_mask) begin
      MEM[MEM_MPORT_3_addr] <= MEM_MPORT_3_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_4_en & MEM_MPORT_4_mask) begin
      MEM[MEM_MPORT_4_addr] <= MEM_MPORT_4_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_5_en & MEM_MPORT_5_mask) begin
      MEM[MEM_MPORT_5_addr] <= MEM_MPORT_5_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_6_en & MEM_MPORT_6_mask) begin
      MEM[MEM_MPORT_6_addr] <= MEM_MPORT_6_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_7_en & MEM_MPORT_7_mask) begin
      MEM[MEM_MPORT_7_addr] <= MEM_MPORT_7_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_8_en & MEM_MPORT_8_mask) begin
      MEM[MEM_MPORT_8_addr] <= MEM_MPORT_8_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_9_en & MEM_MPORT_9_mask) begin
      MEM[MEM_MPORT_9_addr] <= MEM_MPORT_9_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_10_en & MEM_MPORT_10_mask) begin
      MEM[MEM_MPORT_10_addr] <= MEM_MPORT_10_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_11_en & MEM_MPORT_11_mask) begin
      MEM[MEM_MPORT_11_addr] <= MEM_MPORT_11_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_12_en & MEM_MPORT_12_mask) begin
      MEM[MEM_MPORT_12_addr] <= MEM_MPORT_12_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_13_en & MEM_MPORT_13_mask) begin
      MEM[MEM_MPORT_13_addr] <= MEM_MPORT_13_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_14_en & MEM_MPORT_14_mask) begin
      MEM[MEM_MPORT_14_addr] <= MEM_MPORT_14_data; // @[RF.scala 31:15]
    end
    if (MEM_MPORT_15_en & MEM_MPORT_15_mask) begin
      MEM[MEM_MPORT_15_addr] <= MEM_MPORT_15_data; // @[RF.scala 31:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    MEM[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module new_Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input  [63:0] io_in_0_bits_cf_runahead_checkpoint_id,
  input  [4:0]  io_in_0_bits_cf_instrType,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [3:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [2:0]  io_in_0_bits_ctrl_funct3,
  input         io_in_0_bits_ctrl_func24,
  input         io_in_0_bits_ctrl_func23,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc3,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input         io_in_0_bits_ctrl_isMou,
  input  [63:0] io_in_0_bits_data_imm,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_cf_instr,
  input  [38:0] io_in_1_bits_cf_pc,
  input  [38:0] io_in_1_bits_cf_pnpc,
  input         io_in_1_bits_cf_exceptionVec_1,
  input         io_in_1_bits_cf_exceptionVec_2,
  input         io_in_1_bits_cf_exceptionVec_12,
  input         io_in_1_bits_cf_intrVec_0,
  input         io_in_1_bits_cf_intrVec_1,
  input         io_in_1_bits_cf_intrVec_2,
  input         io_in_1_bits_cf_intrVec_3,
  input         io_in_1_bits_cf_intrVec_4,
  input         io_in_1_bits_cf_intrVec_5,
  input         io_in_1_bits_cf_intrVec_6,
  input         io_in_1_bits_cf_intrVec_7,
  input         io_in_1_bits_cf_intrVec_8,
  input         io_in_1_bits_cf_intrVec_9,
  input         io_in_1_bits_cf_intrVec_10,
  input         io_in_1_bits_cf_intrVec_11,
  input  [3:0]  io_in_1_bits_cf_brIdx,
  input         io_in_1_bits_cf_crossPageIPFFix,
  input  [63:0] io_in_1_bits_cf_runahead_checkpoint_id,
  input  [4:0]  io_in_1_bits_cf_instrType,
  input         io_in_1_bits_ctrl_src1Type,
  input         io_in_1_bits_ctrl_src2Type,
  input  [3:0]  io_in_1_bits_ctrl_fuType,
  input  [6:0]  io_in_1_bits_ctrl_fuOpType,
  input  [2:0]  io_in_1_bits_ctrl_funct3,
  input         io_in_1_bits_ctrl_func24,
  input         io_in_1_bits_ctrl_func23,
  input  [4:0]  io_in_1_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_1_bits_ctrl_rfSrc2,
  input  [4:0]  io_in_1_bits_ctrl_rfSrc3,
  input         io_in_1_bits_ctrl_rfWen,
  input  [4:0]  io_in_1_bits_ctrl_rfDest,
  input         io_in_1_bits_ctrl_isMou,
  input  [63:0] io_in_1_bits_data_imm,
  input  [1:0]  io_flush,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  output [1:0]  io_memMMU_imem_priviledgeMode,
  output [1:0]  io_memMMU_dmem_priviledgeMode,
  output        io_memMMU_dmem_status_sum,
  output        io_memMMU_dmem_status_mxr,
  input         io_memMMU_dmem_loadPF,
  input         io_memMMU_dmem_storePF,
  input  [38:0] io_memMMU_dmem_addr,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         _T_408_0,
  output        flushICache,
  output [63:0] perfCnts_2,
  output [38:0] io_in_0_bits_decode_cf_pc,
  output [63:0] satp,
  output        bpuUpdateReq_valid,
  output [38:0] bpuUpdateReq_pc,
  output        bpuUpdateReq_isMissPredict,
  output [38:0] bpuUpdateReq_actualTarget,
  output        bpuUpdateReq_actualTaken,
  output [6:0]  bpuUpdateReq_fuOpType,
  output [1:0]  bpuUpdateReq_btbType,
  output        bpuUpdateReq_isRVC,
  output [4:0]  io_wb_rfDest_0,
  input         ismmio,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  output        io_wb_rfWen_0,
  output [63:0] io_wb_WriteData_0,
  output [63:0] intrVec,
  input         _T_407_0,
  input         io_extra_msip,
  output        flushTLB,
  output        io_in_0_valid_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[Backend.scala 724:20]
  wire  isu_reset; // @[Backend.scala 724:20]
  wire  isu_io_in_0_ready; // @[Backend.scala 724:20]
  wire  isu_io_in_0_valid; // @[Backend.scala 724:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[Backend.scala 724:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[Backend.scala 724:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[Backend.scala 724:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 724:20]
  wire [63:0] isu_io_in_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_0_bits_cf_instrType; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[Backend.scala 724:20]
  wire [3:0] isu_io_in_0_bits_ctrl_fuType; // @[Backend.scala 724:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 724:20]
  wire [2:0] isu_io_in_0_bits_ctrl_funct3; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_ctrl_func24; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_ctrl_func23; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc3; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[Backend.scala 724:20]
  wire  isu_io_in_0_bits_ctrl_isMou; // @[Backend.scala 724:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[Backend.scala 724:20]
  wire  isu_io_in_1_ready; // @[Backend.scala 724:20]
  wire  isu_io_in_1_valid; // @[Backend.scala 724:20]
  wire [63:0] isu_io_in_1_bits_cf_instr; // @[Backend.scala 724:20]
  wire [38:0] isu_io_in_1_bits_cf_pc; // @[Backend.scala 724:20]
  wire [38:0] isu_io_in_1_bits_cf_pnpc; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_exceptionVec_1; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_exceptionVec_2; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_exceptionVec_12; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_0; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_1; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_2; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_3; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_4; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_5; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_6; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_7; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_8; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_9; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_10; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_intrVec_11; // @[Backend.scala 724:20]
  wire [3:0] isu_io_in_1_bits_cf_brIdx; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_cf_crossPageIPFFix; // @[Backend.scala 724:20]
  wire [63:0] isu_io_in_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_1_bits_cf_instrType; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_ctrl_src1Type; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_ctrl_src2Type; // @[Backend.scala 724:20]
  wire [3:0] isu_io_in_1_bits_ctrl_fuType; // @[Backend.scala 724:20]
  wire [6:0] isu_io_in_1_bits_ctrl_fuOpType; // @[Backend.scala 724:20]
  wire [2:0] isu_io_in_1_bits_ctrl_funct3; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_ctrl_func24; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_ctrl_func23; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_1_bits_ctrl_rfSrc1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_1_bits_ctrl_rfSrc2; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_1_bits_ctrl_rfSrc3; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_ctrl_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_in_1_bits_ctrl_rfDest; // @[Backend.scala 724:20]
  wire  isu_io_in_1_bits_ctrl_isMou; // @[Backend.scala 724:20]
  wire [63:0] isu_io_in_1_bits_data_imm; // @[Backend.scala 724:20]
  wire  isu_io_out_0_ready; // @[Backend.scala 724:20]
  wire  isu_io_out_0_valid; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_0_bits_cf_instr; // @[Backend.scala 724:20]
  wire [38:0] isu_io_out_0_bits_cf_pc; // @[Backend.scala 724:20]
  wire [38:0] isu_io_out_0_bits_cf_pnpc; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_exceptionVec_1; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_exceptionVec_2; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_exceptionVec_12; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_0; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_1; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_2; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_3; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_4; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_5; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_6; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_7; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_8; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_9; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_10; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_intrVec_11; // @[Backend.scala 724:20]
  wire [3:0] isu_io_out_0_bits_cf_brIdx; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_cf_crossPageIPFFix; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 724:20]
  wire [4:0] isu_io_out_0_bits_cf_instrType; // @[Backend.scala 724:20]
  wire [3:0] isu_io_out_0_bits_ctrl_fuType; // @[Backend.scala 724:20]
  wire [6:0] isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 724:20]
  wire [2:0] isu_io_out_0_bits_ctrl_funct3; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_ctrl_func24; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_ctrl_func23; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_ctrl_isBru; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_ctrl_isMou; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_0_bits_data_src1; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_0_bits_data_src2; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_0_bits_data_src3; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_0_bits_data_imm; // @[Backend.scala 724:20]
  wire [4:0] isu_io_out_0_bits_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_out_0_bits_InstFlag; // @[Backend.scala 724:20]
  wire  isu_io_out_1_ready; // @[Backend.scala 724:20]
  wire  isu_io_out_1_valid; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_1_bits_cf_instr; // @[Backend.scala 724:20]
  wire [38:0] isu_io_out_1_bits_cf_pc; // @[Backend.scala 724:20]
  wire [38:0] isu_io_out_1_bits_cf_pnpc; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_exceptionVec_1; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_exceptionVec_2; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_exceptionVec_12; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_0; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_1; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_2; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_3; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_4; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_5; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_6; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_7; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_8; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_9; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_10; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_intrVec_11; // @[Backend.scala 724:20]
  wire [3:0] isu_io_out_1_bits_cf_brIdx; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_cf_crossPageIPFFix; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 724:20]
  wire [4:0] isu_io_out_1_bits_cf_instrType; // @[Backend.scala 724:20]
  wire [3:0] isu_io_out_1_bits_ctrl_fuType; // @[Backend.scala 724:20]
  wire [6:0] isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 724:20]
  wire [2:0] isu_io_out_1_bits_ctrl_funct3; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_ctrl_func24; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_ctrl_func23; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_ctrl_isBru; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_ctrl_isMou; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_1_bits_data_src1; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_1_bits_data_src2; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_1_bits_data_src3; // @[Backend.scala 724:20]
  wire [63:0] isu_io_out_1_bits_data_imm; // @[Backend.scala 724:20]
  wire [4:0] isu_io_out_1_bits_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_out_1_bits_InstFlag; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_0; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_1; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_2; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_3; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_4; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_5; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_6; // @[Backend.scala 724:20]
  wire  isu_io_wb_rfWen_7; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_0; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_2; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_3; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_4; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_5; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_6; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfDest_7; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_0; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_1; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_2; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_3; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_4; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_5; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_6; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_WriteData_7; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfSrc1_0; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfSrc1_1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfSrc2_0; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfSrc2_1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfSrc3_0; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_rfSrc3_1; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_ReadData1_0; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_ReadData1_1; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_ReadData2_0; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_ReadData2_1; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_ReadData3_0; // @[Backend.scala 724:20]
  wire [63:0] isu_io_wb_ReadData3_1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_0; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_1; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_2; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_3; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_4; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_5; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_6; // @[Backend.scala 724:20]
  wire [4:0] isu_io_wb_InstNo_7; // @[Backend.scala 724:20]
  wire  isu_io_forward_0_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_0_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_0_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_0_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_0_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_1_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_1_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_1_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_1_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_1_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_2_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_2_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_2_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_2_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_2_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_3_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_3_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_3_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_3_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_3_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_4_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_4_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_4_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_4_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_4_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_5_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_5_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_5_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_5_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_5_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_6_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_6_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_6_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_6_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_6_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_forward_7_valid; // @[Backend.scala 724:20]
  wire  isu_io_forward_7_wb_rfWen; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_7_wb_rfDest; // @[Backend.scala 724:20]
  wire [63:0] isu_io_forward_7_wb_rfData; // @[Backend.scala 724:20]
  wire [4:0] isu_io_forward_7_InstNo; // @[Backend.scala 724:20]
  wire  isu_io_flush; // @[Backend.scala 724:20]
  wire [4:0] isu_io_num_enterwbu; // @[Backend.scala 724:20]
  wire [4:0] isu_io_TailPtr; // @[Backend.scala 724:20]
  wire  exu_clock; // @[Backend.scala 725:20]
  wire  exu_reset; // @[Backend.scala 725:20]
  wire  exu_io__in_0_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_0_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_0_bits_cf_instr; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_0_bits_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_0_bits_cf_pnpc; // @[Backend.scala 725:20]
  wire [3:0] exu_io__in_0_bits_cf_brIdx; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_0_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire  exu_io__in_0_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_0_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_0_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_0_bits_data_src2; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_0_bits_data_imm; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_0_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_0_bits_InstFlag; // @[Backend.scala 725:20]
  wire  exu_io__in_1_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_1_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_1_bits_cf_pc; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_exceptionVec_1; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_exceptionVec_2; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_exceptionVec_12; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_0; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_1; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_2; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_3; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_4; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_5; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_6; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_7; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_8; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_9; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_10; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_intrVec_11; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_cf_crossPageIPFFix; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_1_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_1_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_ctrl_isMou; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_1_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_1_bits_data_src2; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_1_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_1_bits_InstFlag; // @[Backend.scala 725:20]
  wire  exu_io__in_2_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_2_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_2_bits_cf_instr; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_2_bits_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_2_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_2_bits_cf_instrType; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_2_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire [2:0] exu_io__in_2_bits_ctrl_funct3; // @[Backend.scala 725:20]
  wire  exu_io__in_2_bits_ctrl_func24; // @[Backend.scala 725:20]
  wire  exu_io__in_2_bits_ctrl_func23; // @[Backend.scala 725:20]
  wire  exu_io__in_2_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_2_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_2_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_2_bits_data_src2; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_2_bits_data_src3; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_2_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_2_bits_InstFlag; // @[Backend.scala 725:20]
  wire  exu_io__in_3_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_3_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_3_bits_cf_instr; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_3_bits_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_3_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_3_bits_cf_instrType; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_3_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire [2:0] exu_io__in_3_bits_ctrl_funct3; // @[Backend.scala 725:20]
  wire  exu_io__in_3_bits_ctrl_func24; // @[Backend.scala 725:20]
  wire  exu_io__in_3_bits_ctrl_func23; // @[Backend.scala 725:20]
  wire  exu_io__in_3_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_3_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_3_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_3_bits_data_src2; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_3_bits_data_src3; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_3_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_3_bits_InstFlag; // @[Backend.scala 725:20]
  wire  exu_io__in_4_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_4_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_4_bits_cf_instr; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_4_bits_cf_pc; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_exceptionVec_1; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_exceptionVec_2; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_exceptionVec_12; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_0; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_1; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_2; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_3; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_4; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_5; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_6; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_7; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_8; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_9; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_10; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_intrVec_11; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_cf_crossPageIPFFix; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_4_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_4_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_4_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_ctrl_isMou; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_4_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_4_bits_data_src2; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_4_bits_data_imm; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_4_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_4_bits_InstFlag; // @[Backend.scala 725:20]
  wire  exu_io__in_5_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_5_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_5_bits_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_5_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_5_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire  exu_io__in_5_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_5_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_5_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_5_bits_data_src2; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_5_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_6_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_6_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_6_bits_cf_instr; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_6_bits_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_6_bits_cf_pnpc; // @[Backend.scala 725:20]
  wire [3:0] exu_io__in_6_bits_cf_brIdx; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_6_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_6_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire  exu_io__in_6_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_6_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_6_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_6_bits_data_src2; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_6_bits_data_imm; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_6_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__in_7_ready; // @[Backend.scala 725:20]
  wire  exu_io__in_7_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_7_bits_cf_instr; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_7_bits_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__in_7_bits_cf_pnpc; // @[Backend.scala 725:20]
  wire [3:0] exu_io__in_7_bits_cf_brIdx; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_7_bits_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire [6:0] exu_io__in_7_bits_ctrl_fuOpType; // @[Backend.scala 725:20]
  wire  exu_io__in_7_bits_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_7_bits_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_7_bits_data_src1; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_7_bits_data_src2; // @[Backend.scala 725:20]
  wire [63:0] exu_io__in_7_bits_data_imm; // @[Backend.scala 725:20]
  wire [4:0] exu_io__in_7_bits_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__out_0_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_0_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_0_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_0_bits_decode_cf_redirect_target; // @[Backend.scala 725:20]
  wire  exu_io__out_0_bits_decode_cf_redirect_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_0_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_0_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_0_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_0_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__out_0_bits_decode_InstFlag; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_0_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_1_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_1_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_1_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_1_bits_decode_cf_redirect_target; // @[Backend.scala 725:20]
  wire  exu_io__out_1_bits_decode_cf_redirect_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_1_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_1_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_1_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_1_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__out_1_bits_decode_InstFlag; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_1_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_2_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_2_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_2_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_2_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_2_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_2_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire  exu_io__out_2_bits_decode_pext_OV; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_2_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_2_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_3_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_3_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_3_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_3_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_3_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_3_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire  exu_io__out_3_bits_decode_pext_OV; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_3_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_3_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_4_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_4_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_4_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_4_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_4_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_4_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_4_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_4_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_5_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_5_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_5_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_6_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_6_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 725:20]
  wire  exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_6_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__out_7_ready; // @[Backend.scala 725:20]
  wire  exu_io__out_7_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 725:20]
  wire [38:0] exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 725:20]
  wire  exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 725:20]
  wire  exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 725:20]
  wire [4:0] exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 725:20]
  wire [63:0] exu_io__out_7_bits_commits; // @[Backend.scala 725:20]
  wire  exu_io__flush; // @[Backend.scala 725:20]
  wire  exu_io__dmem_req_ready; // @[Backend.scala 725:20]
  wire  exu_io__dmem_req_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[Backend.scala 725:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[Backend.scala 725:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[Backend.scala 725:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[Backend.scala 725:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[Backend.scala 725:20]
  wire  exu_io__dmem_resp_valid; // @[Backend.scala 725:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[Backend.scala 725:20]
  wire  exu_io__forward_0_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_0_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_0_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_0_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_0_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_1_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_1_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_1_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_1_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_1_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_2_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_2_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_2_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_2_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_2_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_3_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_3_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_3_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_3_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_3_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_4_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_4_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_4_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_4_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_4_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_5_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_5_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_5_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_5_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_5_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_6_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_6_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_6_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_6_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_6_InstNo; // @[Backend.scala 725:20]
  wire  exu_io__forward_7_valid; // @[Backend.scala 725:20]
  wire  exu_io__forward_7_wb_rfWen; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_7_wb_rfDest; // @[Backend.scala 725:20]
  wire [63:0] exu_io__forward_7_wb_rfData; // @[Backend.scala 725:20]
  wire [4:0] exu_io__forward_7_InstNo; // @[Backend.scala 725:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 725:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 725:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[Backend.scala 725:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 725:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[Backend.scala 725:20]
  wire  exu_io__memMMU_dmem_storePF; // @[Backend.scala 725:20]
  wire [38:0] exu_io__memMMU_dmem_addr; // @[Backend.scala 725:20]
  wire  exu_lsu_firststage_fire; // @[Backend.scala 725:20]
  wire  exu__T_408; // @[Backend.scala 725:20]
  wire  exu__T_137_0; // @[Backend.scala 725:20]
  wire  exu_flushICache; // @[Backend.scala 725:20]
  wire  exu__T_140_0; // @[Backend.scala 725:20]
  wire [63:0] exu_perfCnts_2; // @[Backend.scala 725:20]
  wire  exu__WIRE_2_0; // @[Backend.scala 725:20]
  wire [63:0] exu_satp; // @[Backend.scala 725:20]
  wire  exu_bpuUpdateReq_valid; // @[Backend.scala 725:20]
  wire [38:0] exu_bpuUpdateReq_pc; // @[Backend.scala 725:20]
  wire  exu_bpuUpdateReq_isMissPredict; // @[Backend.scala 725:20]
  wire [38:0] exu_bpuUpdateReq_actualTarget; // @[Backend.scala 725:20]
  wire  exu_bpuUpdateReq_actualTaken; // @[Backend.scala 725:20]
  wire [6:0] exu_bpuUpdateReq_fuOpType; // @[Backend.scala 725:20]
  wire [1:0] exu_bpuUpdateReq_btbType; // @[Backend.scala 725:20]
  wire  exu_bpuUpdateReq_isRVC; // @[Backend.scala 725:20]
  wire  exu_io_in_0_valid; // @[Backend.scala 725:20]
  wire  exu_ismmio; // @[Backend.scala 725:20]
  wire  exu__WIRE_2_1; // @[Backend.scala 725:20]
  wire  exu_io_extra_mtip; // @[Backend.scala 725:20]
  wire  exu_amoReq; // @[Backend.scala 725:20]
  wire  exu__T_136_0; // @[Backend.scala 725:20]
  wire  exu_io_extra_meip_0; // @[Backend.scala 725:20]
  wire  exu__T_139_0; // @[Backend.scala 725:20]
  wire  exu_vmEnable; // @[Backend.scala 725:20]
  wire [63:0] exu_intrVec; // @[Backend.scala 725:20]
  wire  exu__T_407; // @[Backend.scala 725:20]
  wire  exu__WIRE_1_0; // @[Backend.scala 725:20]
  wire  exu_io_extra_msip; // @[Backend.scala 725:20]
  wire  exu__T_138_0; // @[Backend.scala 725:20]
  wire  exu_flushTLB; // @[Backend.scala 725:20]
  wire  exu__T_135_0; // @[Backend.scala 725:20]
  wire  wbu_clock; // @[Backend.scala 726:20]
  wire  wbu_reset; // @[Backend.scala 726:20]
  wire  wbu_io__in_0_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_0_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_0_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_0_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_0_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_0_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_0_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_0_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_0_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_0_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_1_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_1_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_1_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_1_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_1_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_1_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_1_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_1_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_1_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_1_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_2_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_2_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_2_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_2_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_2_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_2_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_2_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_2_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_2_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_2_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_3_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_3_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_3_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_3_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_3_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_3_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_3_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_3_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_3_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_3_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_4_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_4_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_4_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_4_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_4_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_4_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_4_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_4_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_4_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_4_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_5_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_5_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_5_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_5_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_5_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_5_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_5_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_5_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_5_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_6_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_6_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_6_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_6_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_6_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_6_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_6_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_6_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_6_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__in_7_valid; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_7_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [38:0] wbu_io__in_7_bits_decode_cf_redirect_target; // @[Backend.scala 726:20]
  wire  wbu_io__in_7_bits_decode_cf_redirect_valid; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 726:20]
  wire  wbu_io__in_7_bits_decode_ctrl_rfWen; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_7_bits_decode_ctrl_rfDest; // @[Backend.scala 726:20]
  wire  wbu_io__in_7_bits_decode_pext_OV; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__in_7_bits_decode_InstNo; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__in_7_bits_commits; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_0; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_1; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_2; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_3; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_4; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_5; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_6; // @[Backend.scala 726:20]
  wire  wbu_io__wb_rfWen_7; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_0; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_1; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_2; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_3; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_4; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_5; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_6; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfDest_7; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_0; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_1; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_2; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_3; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_4; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_5; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_6; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_WriteData_7; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfSrc1_0; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfSrc1_1; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfSrc2_0; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfSrc2_1; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfSrc3_0; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_rfSrc3_1; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_ReadData1_0; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_ReadData1_1; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_ReadData2_0; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_ReadData2_1; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_ReadData3_0; // @[Backend.scala 726:20]
  wire [63:0] wbu_io__wb_ReadData3_1; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_0; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_1; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_2; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_3; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_4; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_5; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_6; // @[Backend.scala 726:20]
  wire [4:0] wbu_io__wb_InstNo_7; // @[Backend.scala 726:20]
  wire  wbu_io__redirect_valid; // @[Backend.scala 726:20]
  wire  wbu__T_137_0; // @[Backend.scala 726:20]
  wire  wbu__T_140_0; // @[Backend.scala 726:20]
  wire [38:0] wbu_io_in_0_bits_decode_cf_pc; // @[Backend.scala 726:20]
  wire [4:0] wbu_io_wb_rfDest_0; // @[Backend.scala 726:20]
  wire  wbu_io_in_0_valid; // @[Backend.scala 726:20]
  wire  wbu__WIRE_2_1; // @[Backend.scala 726:20]
  wire  wbu__T_136_0; // @[Backend.scala 726:20]
  wire  wbu__T_139_0; // @[Backend.scala 726:20]
  wire  wbu_io_wb_rfWen_0; // @[Backend.scala 726:20]
  wire [63:0] wbu_io_wb_WriteData_0; // @[Backend.scala 726:20]
  wire  wbu__T_138_0; // @[Backend.scala 726:20]
  wire  wbu_io_in_0_valid_0; // @[Backend.scala 726:20]
  wire  wbu__T_135_0; // @[Backend.scala 726:20]
  reg [63:0] exu_bits_0_cf_instr; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_0_cf_pc; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_0_cf_pnpc; // @[Backend.scala 732:30]
  reg [3:0] exu_bits_0_cf_brIdx; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_0_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_0_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg  exu_bits_0_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_0_ctrl_rfDest; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_0_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_0_data_src2; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_0_data_imm; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_0_InstNo; // @[Backend.scala 732:30]
  reg  exu_bits_0_InstFlag; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_1_cf_pc; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_exceptionVec_1; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_exceptionVec_2; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_exceptionVec_12; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_0; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_1; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_2; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_3; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_4; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_5; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_6; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_7; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_8; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_9; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_10; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_intrVec_11; // @[Backend.scala 732:30]
  reg  exu_bits_1_cf_crossPageIPFFix; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_1_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_1_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg  exu_bits_1_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_1_ctrl_rfDest; // @[Backend.scala 732:30]
  reg  exu_bits_1_ctrl_isMou; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_1_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_1_data_src2; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_1_InstNo; // @[Backend.scala 732:30]
  reg  exu_bits_1_InstFlag; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_2_cf_instr; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_2_cf_pc; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_2_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_2_cf_instrType; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_2_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg [2:0] exu_bits_2_ctrl_funct3; // @[Backend.scala 732:30]
  reg  exu_bits_2_ctrl_func24; // @[Backend.scala 732:30]
  reg  exu_bits_2_ctrl_func23; // @[Backend.scala 732:30]
  reg  exu_bits_2_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_2_ctrl_rfDest; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_2_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_2_data_src2; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_2_data_src3; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_2_InstNo; // @[Backend.scala 732:30]
  reg  exu_bits_2_InstFlag; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_3_cf_instr; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_3_cf_pc; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_3_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_3_cf_instrType; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_3_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg [2:0] exu_bits_3_ctrl_funct3; // @[Backend.scala 732:30]
  reg  exu_bits_3_ctrl_func24; // @[Backend.scala 732:30]
  reg  exu_bits_3_ctrl_func23; // @[Backend.scala 732:30]
  reg  exu_bits_3_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_3_ctrl_rfDest; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_3_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_3_data_src2; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_3_data_src3; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_3_InstNo; // @[Backend.scala 732:30]
  reg  exu_bits_3_InstFlag; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_4_cf_instr; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_4_cf_pc; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_exceptionVec_1; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_exceptionVec_2; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_exceptionVec_12; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_0; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_1; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_2; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_3; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_4; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_5; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_6; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_7; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_8; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_9; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_10; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_intrVec_11; // @[Backend.scala 732:30]
  reg  exu_bits_4_cf_crossPageIPFFix; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_4_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_4_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg  exu_bits_4_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_4_ctrl_rfDest; // @[Backend.scala 732:30]
  reg  exu_bits_4_ctrl_isMou; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_4_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_4_data_src2; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_4_data_imm; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_4_InstNo; // @[Backend.scala 732:30]
  reg  exu_bits_4_InstFlag; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_5_cf_pc; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_5_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_5_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg  exu_bits_5_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_5_ctrl_rfDest; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_5_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_5_data_src2; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_5_InstNo; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_6_cf_instr; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_6_cf_pc; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_6_cf_pnpc; // @[Backend.scala 732:30]
  reg [3:0] exu_bits_6_cf_brIdx; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_6_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_6_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg  exu_bits_6_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_6_ctrl_rfDest; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_6_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_6_data_src2; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_6_data_imm; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_6_InstNo; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_7_cf_instr; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_7_cf_pc; // @[Backend.scala 732:30]
  reg [38:0] exu_bits_7_cf_pnpc; // @[Backend.scala 732:30]
  reg [3:0] exu_bits_7_cf_brIdx; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_7_cf_runahead_checkpoint_id; // @[Backend.scala 732:30]
  reg [6:0] exu_bits_7_ctrl_fuOpType; // @[Backend.scala 732:30]
  reg  exu_bits_7_ctrl_rfWen; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_7_ctrl_rfDest; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_7_data_src1; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_7_data_src2; // @[Backend.scala 732:30]
  reg [63:0] exu_bits_7_data_imm; // @[Backend.scala 732:30]
  reg [4:0] exu_bits_7_InstNo; // @[Backend.scala 732:30]
  reg  exu_valid_0; // @[Backend.scala 734:22]
  reg  exu_valid_1; // @[Backend.scala 734:22]
  reg  exu_valid_2; // @[Backend.scala 734:22]
  reg  exu_valid_3; // @[Backend.scala 734:22]
  reg  exu_valid_4; // @[Backend.scala 734:22]
  reg  exu_valid_5; // @[Backend.scala 734:22]
  reg  exu_valid_6; // @[Backend.scala 734:22]
  reg  exu_valid_7; // @[Backend.scala 734:22]
  wire  _T_7 = exu_io__out_0_ready & exu_io__out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T_7 ? 1'h0 : exu_valid_0; // @[Backend.scala 739:{134,153} 736:50]
  wire  _T_14 = exu_io__out_1_ready & exu_io__out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_14 ? 1'h0 : exu_valid_1; // @[Backend.scala 739:{134,153} 736:50]
  wire  _T_21 = exu_io__out_2_ready & exu_io__out_2_valid; // @[Decoupled.scala 40:37]
  wire  _T_28 = exu_io__out_3_ready & exu_io__out_3_valid; // @[Decoupled.scala 40:37]
  wire  _T_35 = exu_io__out_4_ready & exu_io__out_4_valid; // @[Decoupled.scala 40:37]
  wire  _T_42 = exu_io__out_5_ready & exu_io__out_5_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_42 ? 1'h0 : exu_valid_5; // @[Backend.scala 739:{134,153} 736:50]
  wire  _T_49 = exu_io__out_6_ready & exu_io__out_6_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_49 ? 1'h0 : exu_valid_6; // @[Backend.scala 739:{134,153} 736:50]
  wire  _T_56 = exu_io__out_7_ready & exu_io__out_7_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_56 ? 1'h0 : exu_valid_7; // @[Backend.scala 739:{134,153} 736:50]
  wire  lsu_firststage_fire_0 = exu_lsu_firststage_fire;
  wire  _GEN_8 = lsu_firststage_fire_0 ? 1'h0 : exu_valid_4; // @[Backend.scala 748:{28,56}]
  wire  simdu_fs_fire = exu__WIRE_1_0;
  wire  _GEN_9 = simdu_fs_fire ? 1'h0 : exu_valid_2; // @[Backend.scala 754:{32,62}]
  wire  simdu1_fs_fire = exu__WIRE_2_0;
  wire  _GEN_10 = simdu1_fs_fire ? 1'h0 : exu_valid_3; // @[Backend.scala 757:{35,66}]
  wire  _T_63 = isu_io_out_0_ready & isu_io_out_0_valid; // @[Decoupled.scala 40:37]
  wire  FrontisClear_1 = _T_63 | ~isu_io_in_0_valid; // @[Backend.scala 785:94]
  wire  _T_86 = isu_io_out_0_bits_ctrl_fuType == 4'h6; // @[Backend.scala 762:83]
  wire  _T_93 = isu_io_out_0_bits_ctrl_fuType == 4'h2; // @[Backend.scala 763:84]
  wire  _T_99 = isu_io_out_0_bits_ctrl_fuType == 4'h8; // @[Backend.scala 764:84]
  wire  match_operaotr_0_0 = isu_io_out_0_valid & exu_io__in_0_ready & isu_io_out_0_bits_ctrl_fuType == 4'h0; // @[Backend.scala 805:112]
  wire  match_operaotr_0_1 = ~match_operaotr_0_0 & isu_io_out_0_valid & exu_io__in_1_ready & (
    isu_io_out_0_bits_ctrl_fuType == 4'h1 | _T_99); // @[Backend.scala 805:112]
  wire  _T_182 = match_operaotr_0_0 | match_operaotr_0_1; // @[Backend.scala 801:56]
  wire  match_operaotr_0_2 = ~_T_182 & isu_io_out_0_valid & exu_io__in_2_ready & (_T_93 | _T_93); // @[Backend.scala 805:112]
  wire  _T_236 = match_operaotr_0_0 | match_operaotr_0_1 | match_operaotr_0_2; // @[Backend.scala 801:56]
  wire  match_operaotr_0_3 = ~_T_236 & isu_io_out_0_valid & exu_io__in_3_ready & (isu_io_out_0_bits_ctrl_fuType == 4'h3
     | _T_93); // @[Backend.scala 805:112]
  wire  _T_291 = match_operaotr_0_0 | match_operaotr_0_1 | match_operaotr_0_2 | match_operaotr_0_3; // @[Backend.scala 801:56]
  wire  match_operaotr_0_4 = ~_T_291 & isu_io_out_0_valid & exu_io__in_4_ready & isu_io_out_0_bits_ctrl_fuType == 4'h4; // @[Backend.scala 805:112]
  wire  _T_347 = match_operaotr_0_0 | match_operaotr_0_1 | match_operaotr_0_2 | match_operaotr_0_3 | match_operaotr_0_4; // @[Backend.scala 801:56]
  wire  match_operaotr_0_5 = ~_T_347 & isu_io_out_0_valid & exu_io__in_5_ready & isu_io_out_0_bits_ctrl_fuType == 4'h5; // @[Backend.scala 805:112]
  wire  _T_404 = match_operaotr_0_0 | match_operaotr_0_1 | match_operaotr_0_2 | match_operaotr_0_3 | match_operaotr_0_4
     | match_operaotr_0_5; // @[Backend.scala 801:56]
  wire  _T_419 = isu_io_out_0_bits_ctrl_fuType == 4'h6 & ~isu_io_out_0_bits_ctrl_isBru; // @[Backend.scala 762:153]
  wire  match_operaotr_0_6 = ~_T_404 & isu_io_out_0_valid & exu_io__in_6_ready & (_T_86 | _T_419); // @[Backend.scala 805:112]
  wire  _T_462 = match_operaotr_0_0 | match_operaotr_0_1 | match_operaotr_0_2 | match_operaotr_0_3 | match_operaotr_0_4
     | match_operaotr_0_5 | match_operaotr_0_6; // @[Backend.scala 801:56]
  wire  match_operaotr_0_7 = ~_T_462 & isu_io_out_0_valid & exu_io__in_7_ready & (isu_io_out_0_bits_ctrl_fuType == 4'h7
     | _T_419); // @[Backend.scala 805:112]
  wire  _T_523 = isu_io_out_1_bits_ctrl_fuType == 4'h6; // @[Backend.scala 762:83]
  wire  _T_530 = isu_io_out_1_bits_ctrl_fuType == 4'h2; // @[Backend.scala 763:84]
  wire  _T_536 = isu_io_out_1_bits_ctrl_fuType == 4'h8; // @[Backend.scala 764:84]
  wire  match_operaotr_1_0 = FrontisClear_1 & ~match_operaotr_0_0 & isu_io_out_1_valid & exu_io__in_0_ready &
    isu_io_out_1_bits_ctrl_fuType == 4'h0; // @[Backend.scala 805:112]
  wire  exu_valid_next_0 = match_operaotr_1_0 | (match_operaotr_0_0 | _GEN_0); // @[Backend.scala 805:244 809:29]
  wire  match_operaotr_1_1 = FrontisClear_1 & ~match_operaotr_0_1 & ~match_operaotr_1_0 & isu_io_out_1_valid &
    exu_io__in_1_ready & (isu_io_out_1_bits_ctrl_fuType == 4'h1 | _T_536); // @[Backend.scala 805:112]
  wire  exu_valid_next_1 = match_operaotr_1_1 | (match_operaotr_0_1 | _GEN_1); // @[Backend.scala 805:244 809:29]
  wire  _T_620 = match_operaotr_1_0 | match_operaotr_1_1; // @[Backend.scala 801:56]
  wire  match_operaotr_1_2 = FrontisClear_1 & ~match_operaotr_0_2 & ~_T_620 & isu_io_out_1_valid & exu_io__in_2_ready &
    (_T_530 | _T_530); // @[Backend.scala 805:112]
  wire  exu_valid_next_2 = match_operaotr_1_2 | (match_operaotr_0_2 | _GEN_9); // @[Backend.scala 805:244 809:29]
  wire  _T_675 = match_operaotr_1_0 | match_operaotr_1_1 | match_operaotr_1_2; // @[Backend.scala 801:56]
  wire  match_operaotr_1_3 = FrontisClear_1 & ~match_operaotr_0_3 & ~_T_675 & isu_io_out_1_valid & exu_io__in_3_ready &
    (isu_io_out_1_bits_ctrl_fuType == 4'h3 | _T_530); // @[Backend.scala 805:112]
  wire  exu_valid_next_3 = match_operaotr_1_3 | (match_operaotr_0_3 | _GEN_10); // @[Backend.scala 805:244 809:29]
  wire  _T_731 = match_operaotr_1_0 | match_operaotr_1_1 | match_operaotr_1_2 | match_operaotr_1_3; // @[Backend.scala 801:56]
  wire  match_operaotr_1_4 = FrontisClear_1 & ~match_operaotr_0_4 & ~_T_731 & isu_io_out_1_valid & exu_io__in_4_ready &
    isu_io_out_1_bits_ctrl_fuType == 4'h4; // @[Backend.scala 805:112]
  wire  exu_valid_next_4 = match_operaotr_1_4 | (match_operaotr_0_4 | _GEN_8); // @[Backend.scala 805:244 809:29]
  wire  _T_788 = match_operaotr_1_0 | match_operaotr_1_1 | match_operaotr_1_2 | match_operaotr_1_3 | match_operaotr_1_4; // @[Backend.scala 801:56]
  wire  match_operaotr_1_5 = FrontisClear_1 & ~match_operaotr_0_5 & ~_T_788 & isu_io_out_1_valid & exu_io__in_5_ready &
    isu_io_out_1_bits_ctrl_fuType == 4'h5; // @[Backend.scala 805:112]
  wire  exu_valid_next_5 = match_operaotr_1_5 | (match_operaotr_0_5 | _GEN_5); // @[Backend.scala 805:244 809:29]
  wire  _T_846 = match_operaotr_1_0 | match_operaotr_1_1 | match_operaotr_1_2 | match_operaotr_1_3 | match_operaotr_1_4
     | match_operaotr_1_5; // @[Backend.scala 801:56]
  wire  _T_862 = isu_io_out_1_bits_ctrl_fuType == 4'h6 & ~isu_io_out_1_bits_ctrl_isBru; // @[Backend.scala 762:153]
  wire  match_operaotr_1_6 = FrontisClear_1 & ~match_operaotr_0_6 & ~_T_846 & isu_io_out_1_valid & exu_io__in_6_ready &
    (_T_523 | _T_862); // @[Backend.scala 805:112]
  wire  exu_valid_next_6 = match_operaotr_1_6 | (match_operaotr_0_6 | _GEN_6); // @[Backend.scala 805:244 809:29]
  wire  _T_905 = match_operaotr_1_0 | match_operaotr_1_1 | match_operaotr_1_2 | match_operaotr_1_3 | match_operaotr_1_4
     | match_operaotr_1_5 | match_operaotr_1_6; // @[Backend.scala 801:56]
  wire  match_operaotr_1_7 = FrontisClear_1 & ~match_operaotr_0_7 & ~_T_905 & isu_io_out_1_valid & exu_io__in_7_ready &
    (isu_io_out_1_bits_ctrl_fuType == 4'h7 | _T_862); // @[Backend.scala 805:112]
  wire  exu_valid_next_7 = match_operaotr_1_7 | (match_operaotr_0_7 | _GEN_7); // @[Backend.scala 805:244 809:29]
  wire  _T_964 = exu_io__out_1_bits_decode_InstNo <= exu_io__out_0_bits_decode_InstNo ^
    exu_io__out_1_bits_decode_InstFlag != exu_io__out_0_bits_decode_InstFlag; // @[Backend.scala 826:80]
  wire  _T_966 = exu_io__out_0_valid ? _T_964 : 1'h1; // @[Backend.scala 828:30]
  wire  redirct_index = exu_io__out_1_valid & _T_966; // @[Backend.scala 827:26]
  reg [38:0] wbu_bits_0_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_0_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_0_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_0_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_0_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_0_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_0_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_0_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_0_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_1_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_1_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_1_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_1_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_1_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_1_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_1_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_1_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_1_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_2_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_2_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_2_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_2_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_2_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_2_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_2_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_2_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_2_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_3_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_3_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_3_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_3_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_3_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_3_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_3_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_3_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_3_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_4_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_4_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_4_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_4_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_4_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_4_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_4_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_4_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_4_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_5_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_5_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_5_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_5_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_5_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_5_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_5_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_5_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_5_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_6_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_6_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_6_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_6_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_6_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_6_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_6_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_6_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_6_commits; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_7_decode_cf_pc; // @[Backend.scala 833:30]
  reg [38:0] wbu_bits_7_decode_cf_redirect_target; // @[Backend.scala 833:30]
  reg  wbu_bits_7_decode_cf_redirect_valid; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_7_decode_cf_runahead_checkpoint_id; // @[Backend.scala 833:30]
  reg  wbu_bits_7_decode_ctrl_rfWen; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_7_decode_ctrl_rfDest; // @[Backend.scala 833:30]
  reg  wbu_bits_7_decode_pext_OV; // @[Backend.scala 833:30]
  reg [4:0] wbu_bits_7_decode_InstNo; // @[Backend.scala 833:30]
  reg [63:0] wbu_bits_7_commits; // @[Backend.scala 833:30]
  reg  wbu_valid_0; // @[Backend.scala 835:22]
  reg  wbu_valid_1; // @[Backend.scala 835:22]
  reg  wbu_valid_2; // @[Backend.scala 835:22]
  reg  wbu_valid_3; // @[Backend.scala 835:22]
  reg  wbu_valid_4; // @[Backend.scala 835:22]
  reg  wbu_valid_5; // @[Backend.scala 835:22]
  reg  wbu_valid_6; // @[Backend.scala 835:22]
  reg  wbu_valid_7; // @[Backend.scala 835:22]
  wire [5:0] _GEN_5792 = {{1'd0}, isu_io_TailPtr}; // @[Backend.scala 849:30]
  wire [5:0] ptrleft = 6'h20 - _GEN_5792; // @[Backend.scala 849:30]
  wire [5:0] _GEN_5793 = {{1'd0}, exu_io__out_0_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_973 = _GEN_5793 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_975 = 6'h1 <= ptrleft ? _GEN_5793 == _GEN_5792 : _T_973 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_0 = _T_975 & exu_io__out_0_valid; // @[Backend.scala 866:142]
  wire [63:0] _GEN_1130 = match_exuwbu_0_0 ? exu_io__out_0_bits_commits : wbu_bits_0_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_1134 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_0_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_1135 = match_exuwbu_0_0 ? 1'h0 : wbu_bits_0_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_1147 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_0_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_1148 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_0_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_1161 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_0_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_1193 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_0_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_1195 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_0_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_1197 = match_exuwbu_0_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_0_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire [5:0] _GEN_5795 = {{1'd0}, exu_io__out_1_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_984 = _GEN_5795 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_986 = 6'h1 <= ptrleft ? _GEN_5795 == _GEN_5792 : _T_984 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_1 = _T_986 & exu_io__out_1_valid & ~match_exuwbu_0_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1201 = match_exuwbu_0_1 ? exu_io__out_1_bits_commits : _GEN_1130; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1205 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_1134; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1206 = match_exuwbu_0_1 ? 1'h0 : _GEN_1135; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1218 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_1147; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1219 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_1148; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1232 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_1161; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1264 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_1193; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1266 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_1195; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1268 = match_exuwbu_0_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_1197; // @[Backend.scala 866:202 868:26]
  wire  _T_991 = match_exuwbu_0_0 | match_exuwbu_0_1; // @[Backend.scala 864:57]
  wire [5:0] _GEN_5797 = {{1'd0}, exu_io__out_2_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_996 = _GEN_5797 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_998 = 6'h1 <= ptrleft ? _GEN_5797 == _GEN_5792 : _T_996 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_2 = _T_998 & exu_io__out_2_valid & ~_T_991; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1273 = match_exuwbu_0_2 ? exu_io__out_2_bits_commits : _GEN_1201; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1277 = match_exuwbu_0_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_1205; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1278 = match_exuwbu_0_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_1206; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1290 = match_exuwbu_0_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_1218; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1291 = match_exuwbu_0_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_1219; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1304 = match_exuwbu_0_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_1232; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1336 = match_exuwbu_0_2 ? 1'h0 : _GEN_1264; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1338 = match_exuwbu_0_2 ? 39'h0 : _GEN_1266; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1340 = match_exuwbu_0_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_1268; // @[Backend.scala 866:202 868:26]
  wire  _T_1004 = match_exuwbu_0_0 | match_exuwbu_0_1 | match_exuwbu_0_2; // @[Backend.scala 864:57]
  wire [5:0] _GEN_5799 = {{1'd0}, exu_io__out_3_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_1009 = _GEN_5799 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_1011 = 6'h1 <= ptrleft ? _GEN_5799 == _GEN_5792 : _T_1009 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_3 = _T_1011 & exu_io__out_3_valid & ~_T_1004; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1345 = match_exuwbu_0_3 ? exu_io__out_3_bits_commits : _GEN_1273; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1349 = match_exuwbu_0_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_1277; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1350 = match_exuwbu_0_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_1278; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1362 = match_exuwbu_0_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_1290; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1363 = match_exuwbu_0_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_1291; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1376 = match_exuwbu_0_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_1304; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1408 = match_exuwbu_0_3 ? 1'h0 : _GEN_1336; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1410 = match_exuwbu_0_3 ? 39'h0 : _GEN_1338; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1412 = match_exuwbu_0_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_1340; // @[Backend.scala 866:202 868:26]
  wire  _T_1018 = match_exuwbu_0_0 | match_exuwbu_0_1 | match_exuwbu_0_2 | match_exuwbu_0_3; // @[Backend.scala 864:57]
  wire [5:0] _GEN_5801 = {{1'd0}, exu_io__out_4_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_1023 = _GEN_5801 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_1025 = 6'h1 <= ptrleft ? _GEN_5801 == _GEN_5792 : _T_1023 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_4 = _T_1025 & exu_io__out_4_valid & ~_T_1018; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1417 = match_exuwbu_0_4 ? exu_io__out_4_bits_commits : _GEN_1345; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1421 = match_exuwbu_0_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_1349; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1422 = match_exuwbu_0_4 ? 1'h0 : _GEN_1350; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1434 = match_exuwbu_0_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_1362; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1435 = match_exuwbu_0_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_1363; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1448 = match_exuwbu_0_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_1376; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1480 = match_exuwbu_0_4 ? 1'h0 : _GEN_1408; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1482 = match_exuwbu_0_4 ? 39'h0 : _GEN_1410; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1484 = match_exuwbu_0_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_1412; // @[Backend.scala 866:202 868:26]
  wire  _T_1033 = match_exuwbu_0_0 | match_exuwbu_0_1 | match_exuwbu_0_2 | match_exuwbu_0_3 | match_exuwbu_0_4; // @[Backend.scala 864:57]
  wire [5:0] _GEN_5803 = {{1'd0}, exu_io__out_5_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_1038 = _GEN_5803 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_1040 = 6'h1 <= ptrleft ? _GEN_5803 == _GEN_5792 : _T_1038 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_5 = _T_1040 & exu_io__out_5_valid & ~_T_1033; // @[Backend.scala 866:186]
  wire  _T_1049 = match_exuwbu_0_0 | match_exuwbu_0_1 | match_exuwbu_0_2 | match_exuwbu_0_3 | match_exuwbu_0_4 |
    match_exuwbu_0_5; // @[Backend.scala 864:57]
  wire [5:0] _GEN_5805 = {{1'd0}, exu_io__out_6_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_1054 = _GEN_5805 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_1056 = 6'h1 <= ptrleft ? _GEN_5805 == _GEN_5792 : _T_1054 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_6 = _T_1056 & exu_io__out_6_valid & ~_T_1049; // @[Backend.scala 866:186]
  wire  _T_1066 = match_exuwbu_0_0 | match_exuwbu_0_1 | match_exuwbu_0_2 | match_exuwbu_0_3 | match_exuwbu_0_4 |
    match_exuwbu_0_5 | match_exuwbu_0_6; // @[Backend.scala 864:57]
  wire [5:0] _GEN_5807 = {{1'd0}, exu_io__out_7_bits_decode_InstNo}; // @[Backend.scala 866:68]
  wire [6:0] _T_1071 = _GEN_5807 + ptrleft; // @[Backend.scala 866:122]
  wire  _T_1073 = 6'h1 <= ptrleft ? _GEN_5807 == _GEN_5792 : _T_1071 == 7'h0; // @[Backend.scala 866:15]
  wire  match_exuwbu_0_7 = _T_1073 & exu_io__out_7_valid & ~_T_1066; // @[Backend.scala 866:186]
  wire  wbu_valid_next_0 = match_exuwbu_0_7 | (match_exuwbu_0_6 | (match_exuwbu_0_5 | (match_exuwbu_0_4 | (
    match_exuwbu_0_3 | (match_exuwbu_0_2 | (match_exuwbu_0_1 | match_exuwbu_0_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_1084 = _T_1066 | match_exuwbu_0_7; // @[Backend.scala 865:81]
  wire [5:0] _T_1086 = isu_io_TailPtr + 5'h1; // @[Backend.scala 866:81]
  wire  _T_1090 = 6'h2 <= ptrleft ? _GEN_5793 == _T_1086 : _T_973 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_0 = _T_1090 & exu_io__out_0_valid & _T_1084; // @[Backend.scala 866:165]
  wire [63:0] _GEN_1705 = match_exuwbu_1_0 ? exu_io__out_0_bits_commits : wbu_bits_1_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_1709 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_1_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_1710 = match_exuwbu_1_0 ? 1'h0 : wbu_bits_1_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_1722 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_1_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_1723 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_1_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_1736 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_1_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_1768 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_1_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_1770 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_1_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_1772 = match_exuwbu_1_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_1_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_1108 = 6'h2 <= ptrleft ? _GEN_5795 == _T_1086 : _T_984 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_1 = _T_1108 & exu_io__out_1_valid & _T_1084 & ~match_exuwbu_1_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1777 = match_exuwbu_1_1 ? exu_io__out_1_bits_commits : _GEN_1705; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1781 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_1709; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1782 = match_exuwbu_1_1 ? 1'h0 : _GEN_1710; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1794 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_1722; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1795 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_1723; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1808 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_1736; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1840 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_1768; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1842 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_1770; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1844 = match_exuwbu_1_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_1772; // @[Backend.scala 866:202 868:26]
  wire  _T_1113 = match_exuwbu_1_0 | match_exuwbu_1_1; // @[Backend.scala 864:57]
  wire  _T_1127 = 6'h2 <= ptrleft ? _GEN_5797 == _T_1086 : _T_996 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_2 = _T_1127 & exu_io__out_2_valid & _T_1084 & ~_T_1113; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1849 = match_exuwbu_1_2 ? exu_io__out_2_bits_commits : _GEN_1777; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1853 = match_exuwbu_1_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_1781; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1854 = match_exuwbu_1_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_1782; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1866 = match_exuwbu_1_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_1794; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1867 = match_exuwbu_1_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_1795; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1880 = match_exuwbu_1_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_1808; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1912 = match_exuwbu_1_2 ? 1'h0 : _GEN_1840; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1914 = match_exuwbu_1_2 ? 39'h0 : _GEN_1842; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1916 = match_exuwbu_1_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_1844; // @[Backend.scala 866:202 868:26]
  wire  _T_1133 = match_exuwbu_1_0 | match_exuwbu_1_1 | match_exuwbu_1_2; // @[Backend.scala 864:57]
  wire  _T_1147 = 6'h2 <= ptrleft ? _GEN_5799 == _T_1086 : _T_1009 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_3 = _T_1147 & exu_io__out_3_valid & _T_1084 & ~_T_1133; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1921 = match_exuwbu_1_3 ? exu_io__out_3_bits_commits : _GEN_1849; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1925 = match_exuwbu_1_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_1853; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1926 = match_exuwbu_1_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_1854; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1938 = match_exuwbu_1_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_1866; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1939 = match_exuwbu_1_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_1867; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_1952 = match_exuwbu_1_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_1880; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1984 = match_exuwbu_1_3 ? 1'h0 : _GEN_1912; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1986 = match_exuwbu_1_3 ? 39'h0 : _GEN_1914; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_1988 = match_exuwbu_1_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_1916; // @[Backend.scala 866:202 868:26]
  wire  _T_1154 = match_exuwbu_1_0 | match_exuwbu_1_1 | match_exuwbu_1_2 | match_exuwbu_1_3; // @[Backend.scala 864:57]
  wire  _T_1168 = 6'h2 <= ptrleft ? _GEN_5801 == _T_1086 : _T_1023 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_4 = _T_1168 & exu_io__out_4_valid & _T_1084 & ~_T_1154; // @[Backend.scala 866:186]
  wire [63:0] _GEN_1993 = match_exuwbu_1_4 ? exu_io__out_4_bits_commits : _GEN_1921; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_1997 = match_exuwbu_1_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_1925; // @[Backend.scala 866:202 868:26]
  wire  _GEN_1998 = match_exuwbu_1_4 ? 1'h0 : _GEN_1926; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2010 = match_exuwbu_1_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_1938; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2011 = match_exuwbu_1_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_1939; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_2024 = match_exuwbu_1_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_1952; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2056 = match_exuwbu_1_4 ? 1'h0 : _GEN_1984; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2058 = match_exuwbu_1_4 ? 39'h0 : _GEN_1986; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2060 = match_exuwbu_1_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_1988; // @[Backend.scala 866:202 868:26]
  wire  _T_1176 = match_exuwbu_1_0 | match_exuwbu_1_1 | match_exuwbu_1_2 | match_exuwbu_1_3 | match_exuwbu_1_4; // @[Backend.scala 864:57]
  wire  _T_1190 = 6'h2 <= ptrleft ? _GEN_5803 == _T_1086 : _T_1038 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_5 = _T_1190 & exu_io__out_5_valid & _T_1084 & ~_T_1176; // @[Backend.scala 866:186]
  wire  _T_1199 = match_exuwbu_1_0 | match_exuwbu_1_1 | match_exuwbu_1_2 | match_exuwbu_1_3 | match_exuwbu_1_4 |
    match_exuwbu_1_5; // @[Backend.scala 864:57]
  wire  _T_1213 = 6'h2 <= ptrleft ? _GEN_5805 == _T_1086 : _T_1054 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_6 = _T_1213 & exu_io__out_6_valid & _T_1084 & ~_T_1199; // @[Backend.scala 866:186]
  wire  _T_1223 = match_exuwbu_1_0 | match_exuwbu_1_1 | match_exuwbu_1_2 | match_exuwbu_1_3 | match_exuwbu_1_4 |
    match_exuwbu_1_5 | match_exuwbu_1_6; // @[Backend.scala 864:57]
  wire  _T_1237 = 6'h2 <= ptrleft ? _GEN_5807 == _T_1086 : _T_1071 == 7'h1; // @[Backend.scala 866:15]
  wire  match_exuwbu_1_7 = _T_1237 & exu_io__out_7_valid & _T_1084 & ~_T_1223; // @[Backend.scala 866:186]
  wire  wbu_valid_next_1 = match_exuwbu_1_7 | (match_exuwbu_1_6 | (match_exuwbu_1_5 | (match_exuwbu_1_4 | (
    match_exuwbu_1_3 | (match_exuwbu_1_2 | (match_exuwbu_1_1 | match_exuwbu_1_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_1248 = _T_1223 | match_exuwbu_1_7; // @[Backend.scala 865:81]
  wire [5:0] _T_1250 = isu_io_TailPtr + 5'h2; // @[Backend.scala 866:81]
  wire  _T_1254 = 6'h3 <= ptrleft ? _GEN_5793 == _T_1250 : _T_973 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_0 = _T_1254 & exu_io__out_0_valid & _T_1248; // @[Backend.scala 866:165]
  wire [63:0] _GEN_2281 = match_exuwbu_2_0 ? exu_io__out_0_bits_commits : wbu_bits_2_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_2285 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_2_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_2286 = match_exuwbu_2_0 ? 1'h0 : wbu_bits_2_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_2298 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_2_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_2299 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_2_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_2312 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_2_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_2344 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_2_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_2346 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_2_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_2348 = match_exuwbu_2_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_2_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_1272 = 6'h3 <= ptrleft ? _GEN_5795 == _T_1250 : _T_984 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_1 = _T_1272 & exu_io__out_1_valid & _T_1248 & ~match_exuwbu_2_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_2353 = match_exuwbu_2_1 ? exu_io__out_1_bits_commits : _GEN_2281; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2357 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_2285; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2358 = match_exuwbu_2_1 ? 1'h0 : _GEN_2286; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2370 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_2298; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2371 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_2299; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_2384 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_2312; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2416 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_2344; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2418 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_2346; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2420 = match_exuwbu_2_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_2348; // @[Backend.scala 866:202 868:26]
  wire  _T_1277 = match_exuwbu_2_0 | match_exuwbu_2_1; // @[Backend.scala 864:57]
  wire  _T_1291 = 6'h3 <= ptrleft ? _GEN_5797 == _T_1250 : _T_996 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_2 = _T_1291 & exu_io__out_2_valid & _T_1248 & ~_T_1277; // @[Backend.scala 866:186]
  wire [63:0] _GEN_2425 = match_exuwbu_2_2 ? exu_io__out_2_bits_commits : _GEN_2353; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2429 = match_exuwbu_2_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_2357; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2430 = match_exuwbu_2_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_2358; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2442 = match_exuwbu_2_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_2370; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2443 = match_exuwbu_2_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_2371; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_2456 = match_exuwbu_2_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_2384; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2488 = match_exuwbu_2_2 ? 1'h0 : _GEN_2416; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2490 = match_exuwbu_2_2 ? 39'h0 : _GEN_2418; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2492 = match_exuwbu_2_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_2420; // @[Backend.scala 866:202 868:26]
  wire  _T_1297 = match_exuwbu_2_0 | match_exuwbu_2_1 | match_exuwbu_2_2; // @[Backend.scala 864:57]
  wire  _T_1311 = 6'h3 <= ptrleft ? _GEN_5799 == _T_1250 : _T_1009 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_3 = _T_1311 & exu_io__out_3_valid & _T_1248 & ~_T_1297; // @[Backend.scala 866:186]
  wire [63:0] _GEN_2497 = match_exuwbu_2_3 ? exu_io__out_3_bits_commits : _GEN_2425; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2501 = match_exuwbu_2_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_2429; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2502 = match_exuwbu_2_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_2430; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2514 = match_exuwbu_2_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_2442; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2515 = match_exuwbu_2_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_2443; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_2528 = match_exuwbu_2_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_2456; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2560 = match_exuwbu_2_3 ? 1'h0 : _GEN_2488; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2562 = match_exuwbu_2_3 ? 39'h0 : _GEN_2490; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2564 = match_exuwbu_2_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_2492; // @[Backend.scala 866:202 868:26]
  wire  _T_1318 = match_exuwbu_2_0 | match_exuwbu_2_1 | match_exuwbu_2_2 | match_exuwbu_2_3; // @[Backend.scala 864:57]
  wire  _T_1332 = 6'h3 <= ptrleft ? _GEN_5801 == _T_1250 : _T_1023 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_4 = _T_1332 & exu_io__out_4_valid & _T_1248 & ~_T_1318; // @[Backend.scala 866:186]
  wire [63:0] _GEN_2569 = match_exuwbu_2_4 ? exu_io__out_4_bits_commits : _GEN_2497; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2573 = match_exuwbu_2_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_2501; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2574 = match_exuwbu_2_4 ? 1'h0 : _GEN_2502; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2586 = match_exuwbu_2_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_2514; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2587 = match_exuwbu_2_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_2515; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_2600 = match_exuwbu_2_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_2528; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2632 = match_exuwbu_2_4 ? 1'h0 : _GEN_2560; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2634 = match_exuwbu_2_4 ? 39'h0 : _GEN_2562; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2636 = match_exuwbu_2_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_2564; // @[Backend.scala 866:202 868:26]
  wire  _T_1340 = match_exuwbu_2_0 | match_exuwbu_2_1 | match_exuwbu_2_2 | match_exuwbu_2_3 | match_exuwbu_2_4; // @[Backend.scala 864:57]
  wire  _T_1354 = 6'h3 <= ptrleft ? _GEN_5803 == _T_1250 : _T_1038 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_5 = _T_1354 & exu_io__out_5_valid & _T_1248 & ~_T_1340; // @[Backend.scala 866:186]
  wire  _T_1363 = match_exuwbu_2_0 | match_exuwbu_2_1 | match_exuwbu_2_2 | match_exuwbu_2_3 | match_exuwbu_2_4 |
    match_exuwbu_2_5; // @[Backend.scala 864:57]
  wire  _T_1377 = 6'h3 <= ptrleft ? _GEN_5805 == _T_1250 : _T_1054 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_6 = _T_1377 & exu_io__out_6_valid & _T_1248 & ~_T_1363; // @[Backend.scala 866:186]
  wire  _T_1387 = match_exuwbu_2_0 | match_exuwbu_2_1 | match_exuwbu_2_2 | match_exuwbu_2_3 | match_exuwbu_2_4 |
    match_exuwbu_2_5 | match_exuwbu_2_6; // @[Backend.scala 864:57]
  wire  _T_1401 = 6'h3 <= ptrleft ? _GEN_5807 == _T_1250 : _T_1071 == 7'h2; // @[Backend.scala 866:15]
  wire  match_exuwbu_2_7 = _T_1401 & exu_io__out_7_valid & _T_1248 & ~_T_1387; // @[Backend.scala 866:186]
  wire  wbu_valid_next_2 = match_exuwbu_2_7 | (match_exuwbu_2_6 | (match_exuwbu_2_5 | (match_exuwbu_2_4 | (
    match_exuwbu_2_3 | (match_exuwbu_2_2 | (match_exuwbu_2_1 | match_exuwbu_2_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_1412 = _T_1387 | match_exuwbu_2_7; // @[Backend.scala 865:81]
  wire [5:0] _T_1414 = isu_io_TailPtr + 5'h3; // @[Backend.scala 866:81]
  wire  _T_1418 = 6'h4 <= ptrleft ? _GEN_5793 == _T_1414 : _T_973 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_0 = _T_1418 & exu_io__out_0_valid & _T_1412; // @[Backend.scala 866:165]
  wire [63:0] _GEN_2857 = match_exuwbu_3_0 ? exu_io__out_0_bits_commits : wbu_bits_3_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_2861 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_3_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_2862 = match_exuwbu_3_0 ? 1'h0 : wbu_bits_3_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_2874 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_3_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_2875 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_3_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_2888 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_3_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_2920 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_3_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_2922 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_3_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_2924 = match_exuwbu_3_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_3_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_1436 = 6'h4 <= ptrleft ? _GEN_5795 == _T_1414 : _T_984 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_1 = _T_1436 & exu_io__out_1_valid & _T_1412 & ~match_exuwbu_3_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_2929 = match_exuwbu_3_1 ? exu_io__out_1_bits_commits : _GEN_2857; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2933 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_2861; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2934 = match_exuwbu_3_1 ? 1'h0 : _GEN_2862; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_2946 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_2874; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2947 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_2875; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_2960 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_2888; // @[Backend.scala 866:202 868:26]
  wire  _GEN_2992 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_2920; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2994 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_2922; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_2996 = match_exuwbu_3_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_2924; // @[Backend.scala 866:202 868:26]
  wire  _T_1441 = match_exuwbu_3_0 | match_exuwbu_3_1; // @[Backend.scala 864:57]
  wire  _T_1455 = 6'h4 <= ptrleft ? _GEN_5797 == _T_1414 : _T_996 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_2 = _T_1455 & exu_io__out_2_valid & _T_1412 & ~_T_1441; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3001 = match_exuwbu_3_2 ? exu_io__out_2_bits_commits : _GEN_2929; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3005 = match_exuwbu_3_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_2933; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3006 = match_exuwbu_3_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_2934; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3018 = match_exuwbu_3_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_2946; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3019 = match_exuwbu_3_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_2947; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3032 = match_exuwbu_3_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_2960; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3064 = match_exuwbu_3_2 ? 1'h0 : _GEN_2992; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3066 = match_exuwbu_3_2 ? 39'h0 : _GEN_2994; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3068 = match_exuwbu_3_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_2996; // @[Backend.scala 866:202 868:26]
  wire  _T_1461 = match_exuwbu_3_0 | match_exuwbu_3_1 | match_exuwbu_3_2; // @[Backend.scala 864:57]
  wire  _T_1475 = 6'h4 <= ptrleft ? _GEN_5799 == _T_1414 : _T_1009 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_3 = _T_1475 & exu_io__out_3_valid & _T_1412 & ~_T_1461; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3073 = match_exuwbu_3_3 ? exu_io__out_3_bits_commits : _GEN_3001; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3077 = match_exuwbu_3_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_3005; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3078 = match_exuwbu_3_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_3006; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3090 = match_exuwbu_3_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_3018; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3091 = match_exuwbu_3_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_3019; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3104 = match_exuwbu_3_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_3032; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3136 = match_exuwbu_3_3 ? 1'h0 : _GEN_3064; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3138 = match_exuwbu_3_3 ? 39'h0 : _GEN_3066; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3140 = match_exuwbu_3_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_3068; // @[Backend.scala 866:202 868:26]
  wire  _T_1482 = match_exuwbu_3_0 | match_exuwbu_3_1 | match_exuwbu_3_2 | match_exuwbu_3_3; // @[Backend.scala 864:57]
  wire  _T_1496 = 6'h4 <= ptrleft ? _GEN_5801 == _T_1414 : _T_1023 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_4 = _T_1496 & exu_io__out_4_valid & _T_1412 & ~_T_1482; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3145 = match_exuwbu_3_4 ? exu_io__out_4_bits_commits : _GEN_3073; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3149 = match_exuwbu_3_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_3077; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3150 = match_exuwbu_3_4 ? 1'h0 : _GEN_3078; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3162 = match_exuwbu_3_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_3090; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3163 = match_exuwbu_3_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_3091; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3176 = match_exuwbu_3_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_3104; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3208 = match_exuwbu_3_4 ? 1'h0 : _GEN_3136; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3210 = match_exuwbu_3_4 ? 39'h0 : _GEN_3138; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3212 = match_exuwbu_3_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_3140; // @[Backend.scala 866:202 868:26]
  wire  _T_1504 = match_exuwbu_3_0 | match_exuwbu_3_1 | match_exuwbu_3_2 | match_exuwbu_3_3 | match_exuwbu_3_4; // @[Backend.scala 864:57]
  wire  _T_1518 = 6'h4 <= ptrleft ? _GEN_5803 == _T_1414 : _T_1038 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_5 = _T_1518 & exu_io__out_5_valid & _T_1412 & ~_T_1504; // @[Backend.scala 866:186]
  wire  _T_1527 = match_exuwbu_3_0 | match_exuwbu_3_1 | match_exuwbu_3_2 | match_exuwbu_3_3 | match_exuwbu_3_4 |
    match_exuwbu_3_5; // @[Backend.scala 864:57]
  wire  _T_1541 = 6'h4 <= ptrleft ? _GEN_5805 == _T_1414 : _T_1054 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_6 = _T_1541 & exu_io__out_6_valid & _T_1412 & ~_T_1527; // @[Backend.scala 866:186]
  wire  _T_1551 = match_exuwbu_3_0 | match_exuwbu_3_1 | match_exuwbu_3_2 | match_exuwbu_3_3 | match_exuwbu_3_4 |
    match_exuwbu_3_5 | match_exuwbu_3_6; // @[Backend.scala 864:57]
  wire  _T_1565 = 6'h4 <= ptrleft ? _GEN_5807 == _T_1414 : _T_1071 == 7'h3; // @[Backend.scala 866:15]
  wire  match_exuwbu_3_7 = _T_1565 & exu_io__out_7_valid & _T_1412 & ~_T_1551; // @[Backend.scala 866:186]
  wire  wbu_valid_next_3 = match_exuwbu_3_7 | (match_exuwbu_3_6 | (match_exuwbu_3_5 | (match_exuwbu_3_4 | (
    match_exuwbu_3_3 | (match_exuwbu_3_2 | (match_exuwbu_3_1 | match_exuwbu_3_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_1576 = _T_1551 | match_exuwbu_3_7; // @[Backend.scala 865:81]
  wire [5:0] _T_1578 = isu_io_TailPtr + 5'h4; // @[Backend.scala 866:81]
  wire  _T_1582 = 6'h5 <= ptrleft ? _GEN_5793 == _T_1578 : _T_973 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_0 = _T_1582 & exu_io__out_0_valid & _T_1576; // @[Backend.scala 866:165]
  wire [63:0] _GEN_3433 = match_exuwbu_4_0 ? exu_io__out_0_bits_commits : wbu_bits_4_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_3437 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_4_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_3438 = match_exuwbu_4_0 ? 1'h0 : wbu_bits_4_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_3450 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_4_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_3451 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_4_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_3464 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_4_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_3496 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_4_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_3498 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_4_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_3500 = match_exuwbu_4_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_4_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_1600 = 6'h5 <= ptrleft ? _GEN_5795 == _T_1578 : _T_984 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_1 = _T_1600 & exu_io__out_1_valid & _T_1576 & ~match_exuwbu_4_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3505 = match_exuwbu_4_1 ? exu_io__out_1_bits_commits : _GEN_3433; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3509 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_3437; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3510 = match_exuwbu_4_1 ? 1'h0 : _GEN_3438; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3522 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_3450; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3523 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_3451; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3536 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_3464; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3568 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_3496; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3570 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_3498; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3572 = match_exuwbu_4_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_3500; // @[Backend.scala 866:202 868:26]
  wire  _T_1605 = match_exuwbu_4_0 | match_exuwbu_4_1; // @[Backend.scala 864:57]
  wire  _T_1619 = 6'h5 <= ptrleft ? _GEN_5797 == _T_1578 : _T_996 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_2 = _T_1619 & exu_io__out_2_valid & _T_1576 & ~_T_1605; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3577 = match_exuwbu_4_2 ? exu_io__out_2_bits_commits : _GEN_3505; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3581 = match_exuwbu_4_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_3509; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3582 = match_exuwbu_4_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_3510; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3594 = match_exuwbu_4_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_3522; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3595 = match_exuwbu_4_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_3523; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3608 = match_exuwbu_4_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_3536; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3640 = match_exuwbu_4_2 ? 1'h0 : _GEN_3568; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3642 = match_exuwbu_4_2 ? 39'h0 : _GEN_3570; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3644 = match_exuwbu_4_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_3572; // @[Backend.scala 866:202 868:26]
  wire  _T_1625 = match_exuwbu_4_0 | match_exuwbu_4_1 | match_exuwbu_4_2; // @[Backend.scala 864:57]
  wire  _T_1639 = 6'h5 <= ptrleft ? _GEN_5799 == _T_1578 : _T_1009 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_3 = _T_1639 & exu_io__out_3_valid & _T_1576 & ~_T_1625; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3649 = match_exuwbu_4_3 ? exu_io__out_3_bits_commits : _GEN_3577; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3653 = match_exuwbu_4_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_3581; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3654 = match_exuwbu_4_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_3582; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3666 = match_exuwbu_4_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_3594; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3667 = match_exuwbu_4_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_3595; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3680 = match_exuwbu_4_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_3608; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3712 = match_exuwbu_4_3 ? 1'h0 : _GEN_3640; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3714 = match_exuwbu_4_3 ? 39'h0 : _GEN_3642; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3716 = match_exuwbu_4_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_3644; // @[Backend.scala 866:202 868:26]
  wire  _T_1646 = match_exuwbu_4_0 | match_exuwbu_4_1 | match_exuwbu_4_2 | match_exuwbu_4_3; // @[Backend.scala 864:57]
  wire  _T_1660 = 6'h5 <= ptrleft ? _GEN_5801 == _T_1578 : _T_1023 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_4 = _T_1660 & exu_io__out_4_valid & _T_1576 & ~_T_1646; // @[Backend.scala 866:186]
  wire [63:0] _GEN_3721 = match_exuwbu_4_4 ? exu_io__out_4_bits_commits : _GEN_3649; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3725 = match_exuwbu_4_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_3653; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3726 = match_exuwbu_4_4 ? 1'h0 : _GEN_3654; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_3738 = match_exuwbu_4_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_3666; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3739 = match_exuwbu_4_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_3667; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_3752 = match_exuwbu_4_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_3680; // @[Backend.scala 866:202 868:26]
  wire  _GEN_3784 = match_exuwbu_4_4 ? 1'h0 : _GEN_3712; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3786 = match_exuwbu_4_4 ? 39'h0 : _GEN_3714; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_3788 = match_exuwbu_4_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_3716; // @[Backend.scala 866:202 868:26]
  wire  _T_1668 = match_exuwbu_4_0 | match_exuwbu_4_1 | match_exuwbu_4_2 | match_exuwbu_4_3 | match_exuwbu_4_4; // @[Backend.scala 864:57]
  wire  _T_1682 = 6'h5 <= ptrleft ? _GEN_5803 == _T_1578 : _T_1038 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_5 = _T_1682 & exu_io__out_5_valid & _T_1576 & ~_T_1668; // @[Backend.scala 866:186]
  wire  _T_1691 = match_exuwbu_4_0 | match_exuwbu_4_1 | match_exuwbu_4_2 | match_exuwbu_4_3 | match_exuwbu_4_4 |
    match_exuwbu_4_5; // @[Backend.scala 864:57]
  wire  _T_1705 = 6'h5 <= ptrleft ? _GEN_5805 == _T_1578 : _T_1054 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_6 = _T_1705 & exu_io__out_6_valid & _T_1576 & ~_T_1691; // @[Backend.scala 866:186]
  wire  _T_1715 = match_exuwbu_4_0 | match_exuwbu_4_1 | match_exuwbu_4_2 | match_exuwbu_4_3 | match_exuwbu_4_4 |
    match_exuwbu_4_5 | match_exuwbu_4_6; // @[Backend.scala 864:57]
  wire  _T_1729 = 6'h5 <= ptrleft ? _GEN_5807 == _T_1578 : _T_1071 == 7'h4; // @[Backend.scala 866:15]
  wire  match_exuwbu_4_7 = _T_1729 & exu_io__out_7_valid & _T_1576 & ~_T_1715; // @[Backend.scala 866:186]
  wire  wbu_valid_next_4 = match_exuwbu_4_7 | (match_exuwbu_4_6 | (match_exuwbu_4_5 | (match_exuwbu_4_4 | (
    match_exuwbu_4_3 | (match_exuwbu_4_2 | (match_exuwbu_4_1 | match_exuwbu_4_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_1740 = _T_1715 | match_exuwbu_4_7; // @[Backend.scala 865:81]
  wire [5:0] _T_1742 = isu_io_TailPtr + 5'h5; // @[Backend.scala 866:81]
  wire  _T_1746 = 6'h6 <= ptrleft ? _GEN_5793 == _T_1742 : _T_973 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_0 = _T_1746 & exu_io__out_0_valid & _T_1740; // @[Backend.scala 866:165]
  wire [63:0] _GEN_4009 = match_exuwbu_5_0 ? exu_io__out_0_bits_commits : wbu_bits_5_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_4013 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_5_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_4014 = match_exuwbu_5_0 ? 1'h0 : wbu_bits_5_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_4026 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_5_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_4027 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_5_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_4040 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_5_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_4072 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_5_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_4074 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_5_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_4076 = match_exuwbu_5_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_5_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_1764 = 6'h6 <= ptrleft ? _GEN_5795 == _T_1742 : _T_984 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_1 = _T_1764 & exu_io__out_1_valid & _T_1740 & ~match_exuwbu_5_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4081 = match_exuwbu_5_1 ? exu_io__out_1_bits_commits : _GEN_4009; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4085 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_4013; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4086 = match_exuwbu_5_1 ? 1'h0 : _GEN_4014; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4098 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_4026; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4099 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_4027; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4112 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_4040; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4144 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_4072; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4146 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_4074; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4148 = match_exuwbu_5_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_4076; // @[Backend.scala 866:202 868:26]
  wire  _T_1769 = match_exuwbu_5_0 | match_exuwbu_5_1; // @[Backend.scala 864:57]
  wire  _T_1783 = 6'h6 <= ptrleft ? _GEN_5797 == _T_1742 : _T_996 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_2 = _T_1783 & exu_io__out_2_valid & _T_1740 & ~_T_1769; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4153 = match_exuwbu_5_2 ? exu_io__out_2_bits_commits : _GEN_4081; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4157 = match_exuwbu_5_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_4085; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4158 = match_exuwbu_5_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_4086; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4170 = match_exuwbu_5_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_4098; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4171 = match_exuwbu_5_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_4099; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4184 = match_exuwbu_5_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_4112; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4216 = match_exuwbu_5_2 ? 1'h0 : _GEN_4144; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4218 = match_exuwbu_5_2 ? 39'h0 : _GEN_4146; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4220 = match_exuwbu_5_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_4148; // @[Backend.scala 866:202 868:26]
  wire  _T_1789 = match_exuwbu_5_0 | match_exuwbu_5_1 | match_exuwbu_5_2; // @[Backend.scala 864:57]
  wire  _T_1803 = 6'h6 <= ptrleft ? _GEN_5799 == _T_1742 : _T_1009 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_3 = _T_1803 & exu_io__out_3_valid & _T_1740 & ~_T_1789; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4225 = match_exuwbu_5_3 ? exu_io__out_3_bits_commits : _GEN_4153; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4229 = match_exuwbu_5_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_4157; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4230 = match_exuwbu_5_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_4158; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4242 = match_exuwbu_5_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_4170; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4243 = match_exuwbu_5_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_4171; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4256 = match_exuwbu_5_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_4184; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4288 = match_exuwbu_5_3 ? 1'h0 : _GEN_4216; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4290 = match_exuwbu_5_3 ? 39'h0 : _GEN_4218; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4292 = match_exuwbu_5_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_4220; // @[Backend.scala 866:202 868:26]
  wire  _T_1810 = match_exuwbu_5_0 | match_exuwbu_5_1 | match_exuwbu_5_2 | match_exuwbu_5_3; // @[Backend.scala 864:57]
  wire  _T_1824 = 6'h6 <= ptrleft ? _GEN_5801 == _T_1742 : _T_1023 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_4 = _T_1824 & exu_io__out_4_valid & _T_1740 & ~_T_1810; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4297 = match_exuwbu_5_4 ? exu_io__out_4_bits_commits : _GEN_4225; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4301 = match_exuwbu_5_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_4229; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4302 = match_exuwbu_5_4 ? 1'h0 : _GEN_4230; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4314 = match_exuwbu_5_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_4242; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4315 = match_exuwbu_5_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_4243; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4328 = match_exuwbu_5_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_4256; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4360 = match_exuwbu_5_4 ? 1'h0 : _GEN_4288; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4362 = match_exuwbu_5_4 ? 39'h0 : _GEN_4290; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4364 = match_exuwbu_5_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_4292; // @[Backend.scala 866:202 868:26]
  wire  _T_1832 = match_exuwbu_5_0 | match_exuwbu_5_1 | match_exuwbu_5_2 | match_exuwbu_5_3 | match_exuwbu_5_4; // @[Backend.scala 864:57]
  wire  _T_1846 = 6'h6 <= ptrleft ? _GEN_5803 == _T_1742 : _T_1038 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_5 = _T_1846 & exu_io__out_5_valid & _T_1740 & ~_T_1832; // @[Backend.scala 866:186]
  wire  _T_1855 = match_exuwbu_5_0 | match_exuwbu_5_1 | match_exuwbu_5_2 | match_exuwbu_5_3 | match_exuwbu_5_4 |
    match_exuwbu_5_5; // @[Backend.scala 864:57]
  wire  _T_1869 = 6'h6 <= ptrleft ? _GEN_5805 == _T_1742 : _T_1054 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_6 = _T_1869 & exu_io__out_6_valid & _T_1740 & ~_T_1855; // @[Backend.scala 866:186]
  wire  _T_1879 = match_exuwbu_5_0 | match_exuwbu_5_1 | match_exuwbu_5_2 | match_exuwbu_5_3 | match_exuwbu_5_4 |
    match_exuwbu_5_5 | match_exuwbu_5_6; // @[Backend.scala 864:57]
  wire  _T_1893 = 6'h6 <= ptrleft ? _GEN_5807 == _T_1742 : _T_1071 == 7'h5; // @[Backend.scala 866:15]
  wire  match_exuwbu_5_7 = _T_1893 & exu_io__out_7_valid & _T_1740 & ~_T_1879; // @[Backend.scala 866:186]
  wire  wbu_valid_next_5 = match_exuwbu_5_7 | (match_exuwbu_5_6 | (match_exuwbu_5_5 | (match_exuwbu_5_4 | (
    match_exuwbu_5_3 | (match_exuwbu_5_2 | (match_exuwbu_5_1 | match_exuwbu_5_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_1904 = _T_1879 | match_exuwbu_5_7; // @[Backend.scala 865:81]
  wire [5:0] _T_1906 = isu_io_TailPtr + 5'h6; // @[Backend.scala 866:81]
  wire  _T_1910 = 6'h7 <= ptrleft ? _GEN_5793 == _T_1906 : _T_973 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_0 = _T_1910 & exu_io__out_0_valid & _T_1904; // @[Backend.scala 866:165]
  wire [63:0] _GEN_4585 = match_exuwbu_6_0 ? exu_io__out_0_bits_commits : wbu_bits_6_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_4589 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_6_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_4590 = match_exuwbu_6_0 ? 1'h0 : wbu_bits_6_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_4602 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_6_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_4603 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_6_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_4616 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_6_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_4648 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_6_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_4650 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_6_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_4652 = match_exuwbu_6_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_6_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_1928 = 6'h7 <= ptrleft ? _GEN_5795 == _T_1906 : _T_984 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_1 = _T_1928 & exu_io__out_1_valid & _T_1904 & ~match_exuwbu_6_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4657 = match_exuwbu_6_1 ? exu_io__out_1_bits_commits : _GEN_4585; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4661 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_4589; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4662 = match_exuwbu_6_1 ? 1'h0 : _GEN_4590; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4674 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_4602; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4675 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_4603; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4688 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_4616; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4720 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_4648; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4722 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_4650; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4724 = match_exuwbu_6_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_4652; // @[Backend.scala 866:202 868:26]
  wire  _T_1933 = match_exuwbu_6_0 | match_exuwbu_6_1; // @[Backend.scala 864:57]
  wire  _T_1947 = 6'h7 <= ptrleft ? _GEN_5797 == _T_1906 : _T_996 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_2 = _T_1947 & exu_io__out_2_valid & _T_1904 & ~_T_1933; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4729 = match_exuwbu_6_2 ? exu_io__out_2_bits_commits : _GEN_4657; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4733 = match_exuwbu_6_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_4661; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4734 = match_exuwbu_6_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_4662; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4746 = match_exuwbu_6_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_4674; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4747 = match_exuwbu_6_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_4675; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4760 = match_exuwbu_6_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_4688; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4792 = match_exuwbu_6_2 ? 1'h0 : _GEN_4720; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4794 = match_exuwbu_6_2 ? 39'h0 : _GEN_4722; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4796 = match_exuwbu_6_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_4724; // @[Backend.scala 866:202 868:26]
  wire  _T_1953 = match_exuwbu_6_0 | match_exuwbu_6_1 | match_exuwbu_6_2; // @[Backend.scala 864:57]
  wire  _T_1967 = 6'h7 <= ptrleft ? _GEN_5799 == _T_1906 : _T_1009 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_3 = _T_1967 & exu_io__out_3_valid & _T_1904 & ~_T_1953; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4801 = match_exuwbu_6_3 ? exu_io__out_3_bits_commits : _GEN_4729; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4805 = match_exuwbu_6_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_4733; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4806 = match_exuwbu_6_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_4734; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4818 = match_exuwbu_6_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_4746; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4819 = match_exuwbu_6_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_4747; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4832 = match_exuwbu_6_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_4760; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4864 = match_exuwbu_6_3 ? 1'h0 : _GEN_4792; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4866 = match_exuwbu_6_3 ? 39'h0 : _GEN_4794; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4868 = match_exuwbu_6_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_4796; // @[Backend.scala 866:202 868:26]
  wire  _T_1974 = match_exuwbu_6_0 | match_exuwbu_6_1 | match_exuwbu_6_2 | match_exuwbu_6_3; // @[Backend.scala 864:57]
  wire  _T_1988 = 6'h7 <= ptrleft ? _GEN_5801 == _T_1906 : _T_1023 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_4 = _T_1988 & exu_io__out_4_valid & _T_1904 & ~_T_1974; // @[Backend.scala 866:186]
  wire [63:0] _GEN_4873 = match_exuwbu_6_4 ? exu_io__out_4_bits_commits : _GEN_4801; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4877 = match_exuwbu_6_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_4805; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4878 = match_exuwbu_6_4 ? 1'h0 : _GEN_4806; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_4890 = match_exuwbu_6_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_4818; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4891 = match_exuwbu_6_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_4819; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_4904 = match_exuwbu_6_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_4832; // @[Backend.scala 866:202 868:26]
  wire  _GEN_4936 = match_exuwbu_6_4 ? 1'h0 : _GEN_4864; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4938 = match_exuwbu_6_4 ? 39'h0 : _GEN_4866; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_4940 = match_exuwbu_6_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_4868; // @[Backend.scala 866:202 868:26]
  wire  _T_1996 = match_exuwbu_6_0 | match_exuwbu_6_1 | match_exuwbu_6_2 | match_exuwbu_6_3 | match_exuwbu_6_4; // @[Backend.scala 864:57]
  wire  _T_2010 = 6'h7 <= ptrleft ? _GEN_5803 == _T_1906 : _T_1038 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_5 = _T_2010 & exu_io__out_5_valid & _T_1904 & ~_T_1996; // @[Backend.scala 866:186]
  wire  _T_2019 = match_exuwbu_6_0 | match_exuwbu_6_1 | match_exuwbu_6_2 | match_exuwbu_6_3 | match_exuwbu_6_4 |
    match_exuwbu_6_5; // @[Backend.scala 864:57]
  wire  _T_2033 = 6'h7 <= ptrleft ? _GEN_5805 == _T_1906 : _T_1054 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_6 = _T_2033 & exu_io__out_6_valid & _T_1904 & ~_T_2019; // @[Backend.scala 866:186]
  wire  _T_2043 = match_exuwbu_6_0 | match_exuwbu_6_1 | match_exuwbu_6_2 | match_exuwbu_6_3 | match_exuwbu_6_4 |
    match_exuwbu_6_5 | match_exuwbu_6_6; // @[Backend.scala 864:57]
  wire  _T_2057 = 6'h7 <= ptrleft ? _GEN_5807 == _T_1906 : _T_1071 == 7'h6; // @[Backend.scala 866:15]
  wire  match_exuwbu_6_7 = _T_2057 & exu_io__out_7_valid & _T_1904 & ~_T_2043; // @[Backend.scala 866:186]
  wire  wbu_valid_next_6 = match_exuwbu_6_7 | (match_exuwbu_6_6 | (match_exuwbu_6_5 | (match_exuwbu_6_4 | (
    match_exuwbu_6_3 | (match_exuwbu_6_2 | (match_exuwbu_6_1 | match_exuwbu_6_0)))))); // @[Backend.scala 866:202 869:27]
  wire  _T_2068 = _T_2043 | match_exuwbu_6_7; // @[Backend.scala 865:81]
  wire [5:0] _T_2070 = isu_io_TailPtr + 5'h7; // @[Backend.scala 866:81]
  wire  _T_2074 = 6'h8 <= ptrleft ? _GEN_5793 == _T_2070 : _T_973 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_0 = _T_2074 & exu_io__out_0_valid & _T_2068; // @[Backend.scala 866:165]
  wire [63:0] _GEN_5161 = match_exuwbu_7_0 ? exu_io__out_0_bits_commits : wbu_bits_7_commits; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_5165 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_InstNo : wbu_bits_7_decode_InstNo; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_5166 = match_exuwbu_7_0 ? 1'h0 : wbu_bits_7_decode_pext_OV; // @[Backend.scala 834:17 866:202 868:26]
  wire [4:0] _GEN_5178 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_ctrl_rfDest : wbu_bits_7_decode_ctrl_rfDest; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_5179 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_ctrl_rfWen : wbu_bits_7_decode_ctrl_rfWen; // @[Backend.scala 834:17 866:202 868:26]
  wire [63:0] _GEN_5192 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_cf_runahead_checkpoint_id :
    wbu_bits_7_decode_cf_runahead_checkpoint_id; // @[Backend.scala 834:17 866:202 868:26]
  wire  _GEN_5224 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_cf_redirect_valid : wbu_bits_7_decode_cf_redirect_valid
    ; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_5226 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_cf_redirect_target :
    wbu_bits_7_decode_cf_redirect_target; // @[Backend.scala 834:17 866:202 868:26]
  wire [38:0] _GEN_5228 = match_exuwbu_7_0 ? exu_io__out_0_bits_decode_cf_pc : wbu_bits_7_decode_cf_pc; // @[Backend.scala 834:17 866:202 868:26]
  wire  _T_2092 = 6'h8 <= ptrleft ? _GEN_5795 == _T_2070 : _T_984 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_1 = _T_2092 & exu_io__out_1_valid & _T_2068 & ~match_exuwbu_7_0; // @[Backend.scala 866:186]
  wire [63:0] _GEN_5233 = match_exuwbu_7_1 ? exu_io__out_1_bits_commits : _GEN_5161; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5237 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_InstNo : _GEN_5165; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5238 = match_exuwbu_7_1 ? 1'h0 : _GEN_5166; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5250 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_ctrl_rfDest : _GEN_5178; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5251 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_ctrl_rfWen : _GEN_5179; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_5264 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_cf_runahead_checkpoint_id : _GEN_5192; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5296 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_cf_redirect_valid : _GEN_5224; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5298 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_5226; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5300 = match_exuwbu_7_1 ? exu_io__out_1_bits_decode_cf_pc : _GEN_5228; // @[Backend.scala 866:202 868:26]
  wire  _T_2097 = match_exuwbu_7_0 | match_exuwbu_7_1; // @[Backend.scala 864:57]
  wire  _T_2111 = 6'h8 <= ptrleft ? _GEN_5797 == _T_2070 : _T_996 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_2 = _T_2111 & exu_io__out_2_valid & _T_2068 & ~_T_2097; // @[Backend.scala 866:186]
  wire [63:0] _GEN_5305 = match_exuwbu_7_2 ? exu_io__out_2_bits_commits : _GEN_5233; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5309 = match_exuwbu_7_2 ? exu_io__out_2_bits_decode_InstNo : _GEN_5237; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5310 = match_exuwbu_7_2 ? exu_io__out_2_bits_decode_pext_OV : _GEN_5238; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5322 = match_exuwbu_7_2 ? exu_io__out_2_bits_decode_ctrl_rfDest : _GEN_5250; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5323 = match_exuwbu_7_2 ? exu_io__out_2_bits_decode_ctrl_rfWen : _GEN_5251; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_5336 = match_exuwbu_7_2 ? exu_io__out_2_bits_decode_cf_runahead_checkpoint_id : _GEN_5264; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5368 = match_exuwbu_7_2 ? 1'h0 : _GEN_5296; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5370 = match_exuwbu_7_2 ? 39'h0 : _GEN_5298; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5372 = match_exuwbu_7_2 ? exu_io__out_2_bits_decode_cf_pc : _GEN_5300; // @[Backend.scala 866:202 868:26]
  wire  _T_2117 = match_exuwbu_7_0 | match_exuwbu_7_1 | match_exuwbu_7_2; // @[Backend.scala 864:57]
  wire  _T_2131 = 6'h8 <= ptrleft ? _GEN_5799 == _T_2070 : _T_1009 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_3 = _T_2131 & exu_io__out_3_valid & _T_2068 & ~_T_2117; // @[Backend.scala 866:186]
  wire [63:0] _GEN_5377 = match_exuwbu_7_3 ? exu_io__out_3_bits_commits : _GEN_5305; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5381 = match_exuwbu_7_3 ? exu_io__out_3_bits_decode_InstNo : _GEN_5309; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5382 = match_exuwbu_7_3 ? exu_io__out_3_bits_decode_pext_OV : _GEN_5310; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5394 = match_exuwbu_7_3 ? exu_io__out_3_bits_decode_ctrl_rfDest : _GEN_5322; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5395 = match_exuwbu_7_3 ? exu_io__out_3_bits_decode_ctrl_rfWen : _GEN_5323; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_5408 = match_exuwbu_7_3 ? exu_io__out_3_bits_decode_cf_runahead_checkpoint_id : _GEN_5336; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5440 = match_exuwbu_7_3 ? 1'h0 : _GEN_5368; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5442 = match_exuwbu_7_3 ? 39'h0 : _GEN_5370; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5444 = match_exuwbu_7_3 ? exu_io__out_3_bits_decode_cf_pc : _GEN_5372; // @[Backend.scala 866:202 868:26]
  wire  _T_2138 = match_exuwbu_7_0 | match_exuwbu_7_1 | match_exuwbu_7_2 | match_exuwbu_7_3; // @[Backend.scala 864:57]
  wire  _T_2152 = 6'h8 <= ptrleft ? _GEN_5801 == _T_2070 : _T_1023 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_4 = _T_2152 & exu_io__out_4_valid & _T_2068 & ~_T_2138; // @[Backend.scala 866:186]
  wire [63:0] _GEN_5449 = match_exuwbu_7_4 ? exu_io__out_4_bits_commits : _GEN_5377; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5453 = match_exuwbu_7_4 ? exu_io__out_4_bits_decode_InstNo : _GEN_5381; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5454 = match_exuwbu_7_4 ? 1'h0 : _GEN_5382; // @[Backend.scala 866:202 868:26]
  wire [4:0] _GEN_5466 = match_exuwbu_7_4 ? exu_io__out_4_bits_decode_ctrl_rfDest : _GEN_5394; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5467 = match_exuwbu_7_4 ? exu_io__out_4_bits_decode_ctrl_rfWen : _GEN_5395; // @[Backend.scala 866:202 868:26]
  wire [63:0] _GEN_5480 = match_exuwbu_7_4 ? exu_io__out_4_bits_decode_cf_runahead_checkpoint_id : _GEN_5408; // @[Backend.scala 866:202 868:26]
  wire  _GEN_5512 = match_exuwbu_7_4 ? 1'h0 : _GEN_5440; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5514 = match_exuwbu_7_4 ? 39'h0 : _GEN_5442; // @[Backend.scala 866:202 868:26]
  wire [38:0] _GEN_5516 = match_exuwbu_7_4 ? exu_io__out_4_bits_decode_cf_pc : _GEN_5444; // @[Backend.scala 866:202 868:26]
  wire  _T_2160 = match_exuwbu_7_0 | match_exuwbu_7_1 | match_exuwbu_7_2 | match_exuwbu_7_3 | match_exuwbu_7_4; // @[Backend.scala 864:57]
  wire  _T_2174 = 6'h8 <= ptrleft ? _GEN_5803 == _T_2070 : _T_1038 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_5 = _T_2174 & exu_io__out_5_valid & _T_2068 & ~_T_2160; // @[Backend.scala 866:186]
  wire  _T_2183 = match_exuwbu_7_0 | match_exuwbu_7_1 | match_exuwbu_7_2 | match_exuwbu_7_3 | match_exuwbu_7_4 |
    match_exuwbu_7_5; // @[Backend.scala 864:57]
  wire  _T_2197 = 6'h8 <= ptrleft ? _GEN_5805 == _T_2070 : _T_1054 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_6 = _T_2197 & exu_io__out_6_valid & _T_2068 & ~_T_2183; // @[Backend.scala 866:186]
  wire  _T_2207 = match_exuwbu_7_0 | match_exuwbu_7_1 | match_exuwbu_7_2 | match_exuwbu_7_3 | match_exuwbu_7_4 |
    match_exuwbu_7_5 | match_exuwbu_7_6; // @[Backend.scala 864:57]
  wire  _T_2221 = 6'h8 <= ptrleft ? _GEN_5807 == _T_2070 : _T_1071 == 7'h7; // @[Backend.scala 866:15]
  wire  match_exuwbu_7_7 = _T_2221 & exu_io__out_7_valid & _T_2068 & ~_T_2207; // @[Backend.scala 866:186]
  wire  wbu_valid_next_7 = match_exuwbu_7_7 | (match_exuwbu_7_6 | (match_exuwbu_7_5 | (match_exuwbu_7_4 | (
    match_exuwbu_7_3 | (match_exuwbu_7_2 | (match_exuwbu_7_1 | match_exuwbu_7_0)))))); // @[Backend.scala 866:202 869:27]
  wire [4:0] _T_2228 = exu_io__out_4_bits_decode_InstNo - isu_io_TailPtr; // @[Backend.scala 876:119]
  wire [5:0] _T_2230 = _GEN_5801 + ptrleft; // @[Backend.scala 876:171]
  wire [5:0] lsuInstNo = exu_io__out_4_bits_decode_InstNo >= isu_io_TailPtr ? {{1'd0}, _T_2228} : _T_2230; // @[Backend.scala 876:22]
  wire  _GEN_5736 = 6'h0 < lsuInstNo & ~wbu_valid_next_0 ? 1'h0 : 1'h1; // @[Backend.scala 878:48 879:19]
  wire  _GEN_5737 = 6'h1 < lsuInstNo & ~wbu_valid_next_1 ? 1'h0 : _GEN_5736; // @[Backend.scala 878:48 879:19]
  wire  _GEN_5738 = 6'h2 < lsuInstNo & ~wbu_valid_next_2 ? 1'h0 : _GEN_5737; // @[Backend.scala 878:48 879:19]
  wire  _GEN_5739 = 6'h3 < lsuInstNo & ~wbu_valid_next_3 ? 1'h0 : _GEN_5738; // @[Backend.scala 878:48 879:19]
  wire  _GEN_5740 = 6'h4 < lsuInstNo & ~wbu_valid_next_4 ? 1'h0 : _GEN_5739; // @[Backend.scala 878:48 879:19]
  wire  _GEN_5741 = 6'h5 < lsuInstNo & ~wbu_valid_next_5 ? 1'h0 : _GEN_5740; // @[Backend.scala 878:48 879:19]
  wire  _GEN_5742 = 6'h6 < lsuInstNo & ~wbu_valid_next_6 ? 1'h0 : _GEN_5741; // @[Backend.scala 878:48 879:19]
  wire [1:0] _T_2263 = _T_7 + _T_14; // @[Backend.scala 884:67]
  wire [1:0] _GEN_5922 = {{1'd0}, _T_21}; // @[Backend.scala 884:67]
  wire [2:0] _T_2264 = _T_2263 + _GEN_5922; // @[Backend.scala 884:67]
  wire [2:0] _GEN_5923 = {{2'd0}, _T_28}; // @[Backend.scala 884:67]
  wire [3:0] _T_2265 = _T_2264 + _GEN_5923; // @[Backend.scala 884:67]
  wire [3:0] _GEN_5924 = {{3'd0}, _T_35}; // @[Backend.scala 884:67]
  wire [4:0] _T_2266 = _T_2265 + _GEN_5924; // @[Backend.scala 884:67]
  wire [4:0] _GEN_5925 = {{4'd0}, _T_42}; // @[Backend.scala 884:67]
  wire [5:0] _T_2267 = _T_2266 + _GEN_5925; // @[Backend.scala 884:67]
  wire [5:0] _GEN_5926 = {{5'd0}, _T_49}; // @[Backend.scala 884:67]
  wire [6:0] _T_2268 = _T_2267 + _GEN_5926; // @[Backend.scala 884:67]
  wire [6:0] _GEN_5927 = {{6'd0}, _T_56}; // @[Backend.scala 884:67]
  wire [7:0] num_enterwbu = _T_2268 + _GEN_5927; // @[Backend.scala 884:67]
  wire  _GEN_5753 = redirct_index ? exu_io__out_1_bits_decode_cf_redirect_valid :
    exu_io__out_0_bits_decode_cf_redirect_valid; // @[]
  wire [1:0] _GEN_5928 = {{1'd0}, redirct_index}; // @[]
  wire  _GEN_5754 = 2'h2 == _GEN_5928 ? 1'h0 : _GEN_5753; // @[]
  wire  _GEN_5755 = 2'h3 == _GEN_5928 ? 1'h0 : _GEN_5754; // @[]
  wire [2:0] _GEN_5930 = {{2'd0}, redirct_index}; // @[]
  wire  _GEN_5756 = 3'h4 == _GEN_5930 ? 1'h0 : _GEN_5755; // @[]
  wire  _GEN_5757 = 3'h5 == _GEN_5930 ? 1'h0 : _GEN_5756; // @[]
  wire  _GEN_5758 = 3'h6 == _GEN_5930 ? exu_io__out_6_bits_decode_cf_redirect_valid : _GEN_5757; // @[]
  wire  _GEN_5759 = 3'h7 == _GEN_5930 ? exu_io__out_7_bits_decode_cf_redirect_valid : _GEN_5758; // @[]
  wire [38:0] _GEN_5768 = exu_io__out_0_bits_decode_cf_redirect_target; // @[]
  wire [38:0] _GEN_5769 = redirct_index ? exu_io__out_1_bits_decode_cf_redirect_target : _GEN_5768; // @[]
  wire [38:0] _GEN_5770 = 2'h2 == _GEN_5928 ? 39'h0 : _GEN_5769; // @[]
  wire [38:0] _GEN_5771 = 2'h3 == _GEN_5928 ? 39'h0 : _GEN_5770; // @[]
  wire [38:0] _GEN_5772 = 3'h4 == _GEN_5930 ? 39'h0 : _GEN_5771; // @[]
  wire [38:0] _GEN_5773 = 3'h5 == _GEN_5930 ? 39'h0 : _GEN_5772; // @[]
  wire [38:0] _GEN_5774 = 3'h6 == _GEN_5930 ? exu_io__out_6_bits_decode_cf_redirect_target : _GEN_5773; // @[]
  wire  _GEN_5777 = redirct_index ? exu_io__out_1_ready : exu_io__out_0_ready; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5778 = 2'h2 == _GEN_5928 ? exu_io__out_2_ready : _GEN_5777; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5779 = 2'h3 == _GEN_5928 ? exu_io__out_3_ready : _GEN_5778; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5780 = 3'h4 == _GEN_5930 ? exu_io__out_4_ready : _GEN_5779; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5781 = 3'h5 == _GEN_5930 ? exu_io__out_5_ready : _GEN_5780; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5782 = 3'h6 == _GEN_5930 ? exu_io__out_6_ready : _GEN_5781; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5783 = 3'h7 == _GEN_5930 ? exu_io__out_7_ready : _GEN_5782; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5785 = redirct_index ? exu_io__out_1_valid : exu_io__out_0_valid; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5786 = 2'h2 == _GEN_5928 ? exu_io__out_2_valid : _GEN_5785; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5787 = 2'h3 == _GEN_5928 ? exu_io__out_3_valid : _GEN_5786; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5788 = 3'h4 == _GEN_5930 ? exu_io__out_4_valid : _GEN_5787; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5789 = 3'h5 == _GEN_5930 ? exu_io__out_5_valid : _GEN_5788; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5790 = 3'h6 == _GEN_5930 ? exu_io__out_6_valid : _GEN_5789; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5791 = 3'h7 == _GEN_5930 ? exu_io__out_7_valid : _GEN_5790; // @[Decoupled.scala 40:{37,37}]
  wire  _T_2274 = _GEN_5783 & _GEN_5791; // @[Decoupled.scala 40:37]
  new_SIMD_ISU isu ( // @[Backend.scala 724:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(isu_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_cf_runahead_checkpoint_id(isu_io_in_0_bits_cf_runahead_checkpoint_id),
    .io_in_0_bits_cf_instrType(isu_io_in_0_bits_cf_instrType),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_funct3(isu_io_in_0_bits_ctrl_funct3),
    .io_in_0_bits_ctrl_func24(isu_io_in_0_bits_ctrl_func24),
    .io_in_0_bits_ctrl_func23(isu_io_in_0_bits_ctrl_func23),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfSrc3(isu_io_in_0_bits_ctrl_rfSrc3),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isMou(isu_io_in_0_bits_ctrl_isMou),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_in_1_ready(isu_io_in_1_ready),
    .io_in_1_valid(isu_io_in_1_valid),
    .io_in_1_bits_cf_instr(isu_io_in_1_bits_cf_instr),
    .io_in_1_bits_cf_pc(isu_io_in_1_bits_cf_pc),
    .io_in_1_bits_cf_pnpc(isu_io_in_1_bits_cf_pnpc),
    .io_in_1_bits_cf_exceptionVec_1(isu_io_in_1_bits_cf_exceptionVec_1),
    .io_in_1_bits_cf_exceptionVec_2(isu_io_in_1_bits_cf_exceptionVec_2),
    .io_in_1_bits_cf_exceptionVec_12(isu_io_in_1_bits_cf_exceptionVec_12),
    .io_in_1_bits_cf_intrVec_0(isu_io_in_1_bits_cf_intrVec_0),
    .io_in_1_bits_cf_intrVec_1(isu_io_in_1_bits_cf_intrVec_1),
    .io_in_1_bits_cf_intrVec_2(isu_io_in_1_bits_cf_intrVec_2),
    .io_in_1_bits_cf_intrVec_3(isu_io_in_1_bits_cf_intrVec_3),
    .io_in_1_bits_cf_intrVec_4(isu_io_in_1_bits_cf_intrVec_4),
    .io_in_1_bits_cf_intrVec_5(isu_io_in_1_bits_cf_intrVec_5),
    .io_in_1_bits_cf_intrVec_6(isu_io_in_1_bits_cf_intrVec_6),
    .io_in_1_bits_cf_intrVec_7(isu_io_in_1_bits_cf_intrVec_7),
    .io_in_1_bits_cf_intrVec_8(isu_io_in_1_bits_cf_intrVec_8),
    .io_in_1_bits_cf_intrVec_9(isu_io_in_1_bits_cf_intrVec_9),
    .io_in_1_bits_cf_intrVec_10(isu_io_in_1_bits_cf_intrVec_10),
    .io_in_1_bits_cf_intrVec_11(isu_io_in_1_bits_cf_intrVec_11),
    .io_in_1_bits_cf_brIdx(isu_io_in_1_bits_cf_brIdx),
    .io_in_1_bits_cf_crossPageIPFFix(isu_io_in_1_bits_cf_crossPageIPFFix),
    .io_in_1_bits_cf_runahead_checkpoint_id(isu_io_in_1_bits_cf_runahead_checkpoint_id),
    .io_in_1_bits_cf_instrType(isu_io_in_1_bits_cf_instrType),
    .io_in_1_bits_ctrl_src1Type(isu_io_in_1_bits_ctrl_src1Type),
    .io_in_1_bits_ctrl_src2Type(isu_io_in_1_bits_ctrl_src2Type),
    .io_in_1_bits_ctrl_fuType(isu_io_in_1_bits_ctrl_fuType),
    .io_in_1_bits_ctrl_fuOpType(isu_io_in_1_bits_ctrl_fuOpType),
    .io_in_1_bits_ctrl_funct3(isu_io_in_1_bits_ctrl_funct3),
    .io_in_1_bits_ctrl_func24(isu_io_in_1_bits_ctrl_func24),
    .io_in_1_bits_ctrl_func23(isu_io_in_1_bits_ctrl_func23),
    .io_in_1_bits_ctrl_rfSrc1(isu_io_in_1_bits_ctrl_rfSrc1),
    .io_in_1_bits_ctrl_rfSrc2(isu_io_in_1_bits_ctrl_rfSrc2),
    .io_in_1_bits_ctrl_rfSrc3(isu_io_in_1_bits_ctrl_rfSrc3),
    .io_in_1_bits_ctrl_rfWen(isu_io_in_1_bits_ctrl_rfWen),
    .io_in_1_bits_ctrl_rfDest(isu_io_in_1_bits_ctrl_rfDest),
    .io_in_1_bits_ctrl_isMou(isu_io_in_1_bits_ctrl_isMou),
    .io_in_1_bits_data_imm(isu_io_in_1_bits_data_imm),
    .io_out_0_ready(isu_io_out_0_ready),
    .io_out_0_valid(isu_io_out_0_valid),
    .io_out_0_bits_cf_instr(isu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(isu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(isu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(isu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(isu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(isu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(isu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(isu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(isu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(isu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(isu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(isu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(isu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(isu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(isu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(isu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(isu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(isu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(isu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(isu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_runahead_checkpoint_id(isu_io_out_0_bits_cf_runahead_checkpoint_id),
    .io_out_0_bits_cf_instrType(isu_io_out_0_bits_cf_instrType),
    .io_out_0_bits_ctrl_fuType(isu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(isu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_funct3(isu_io_out_0_bits_ctrl_funct3),
    .io_out_0_bits_ctrl_func24(isu_io_out_0_bits_ctrl_func24),
    .io_out_0_bits_ctrl_func23(isu_io_out_0_bits_ctrl_func23),
    .io_out_0_bits_ctrl_rfWen(isu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(isu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isBru(isu_io_out_0_bits_ctrl_isBru),
    .io_out_0_bits_ctrl_isMou(isu_io_out_0_bits_ctrl_isMou),
    .io_out_0_bits_data_src1(isu_io_out_0_bits_data_src1),
    .io_out_0_bits_data_src2(isu_io_out_0_bits_data_src2),
    .io_out_0_bits_data_src3(isu_io_out_0_bits_data_src3),
    .io_out_0_bits_data_imm(isu_io_out_0_bits_data_imm),
    .io_out_0_bits_InstNo(isu_io_out_0_bits_InstNo),
    .io_out_0_bits_InstFlag(isu_io_out_0_bits_InstFlag),
    .io_out_1_ready(isu_io_out_1_ready),
    .io_out_1_valid(isu_io_out_1_valid),
    .io_out_1_bits_cf_instr(isu_io_out_1_bits_cf_instr),
    .io_out_1_bits_cf_pc(isu_io_out_1_bits_cf_pc),
    .io_out_1_bits_cf_pnpc(isu_io_out_1_bits_cf_pnpc),
    .io_out_1_bits_cf_exceptionVec_1(isu_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(isu_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(isu_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_intrVec_0(isu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(isu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(isu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(isu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(isu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(isu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(isu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(isu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(isu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(isu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(isu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(isu_io_out_1_bits_cf_intrVec_11),
    .io_out_1_bits_cf_brIdx(isu_io_out_1_bits_cf_brIdx),
    .io_out_1_bits_cf_crossPageIPFFix(isu_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_cf_runahead_checkpoint_id(isu_io_out_1_bits_cf_runahead_checkpoint_id),
    .io_out_1_bits_cf_instrType(isu_io_out_1_bits_cf_instrType),
    .io_out_1_bits_ctrl_fuType(isu_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(isu_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_funct3(isu_io_out_1_bits_ctrl_funct3),
    .io_out_1_bits_ctrl_func24(isu_io_out_1_bits_ctrl_func24),
    .io_out_1_bits_ctrl_func23(isu_io_out_1_bits_ctrl_func23),
    .io_out_1_bits_ctrl_rfWen(isu_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_rfDest(isu_io_out_1_bits_ctrl_rfDest),
    .io_out_1_bits_ctrl_isBru(isu_io_out_1_bits_ctrl_isBru),
    .io_out_1_bits_ctrl_isMou(isu_io_out_1_bits_ctrl_isMou),
    .io_out_1_bits_data_src1(isu_io_out_1_bits_data_src1),
    .io_out_1_bits_data_src2(isu_io_out_1_bits_data_src2),
    .io_out_1_bits_data_src3(isu_io_out_1_bits_data_src3),
    .io_out_1_bits_data_imm(isu_io_out_1_bits_data_imm),
    .io_out_1_bits_InstNo(isu_io_out_1_bits_InstNo),
    .io_out_1_bits_InstFlag(isu_io_out_1_bits_InstFlag),
    .io_wb_rfWen_0(isu_io_wb_rfWen_0),
    .io_wb_rfWen_1(isu_io_wb_rfWen_1),
    .io_wb_rfWen_2(isu_io_wb_rfWen_2),
    .io_wb_rfWen_3(isu_io_wb_rfWen_3),
    .io_wb_rfWen_4(isu_io_wb_rfWen_4),
    .io_wb_rfWen_5(isu_io_wb_rfWen_5),
    .io_wb_rfWen_6(isu_io_wb_rfWen_6),
    .io_wb_rfWen_7(isu_io_wb_rfWen_7),
    .io_wb_rfDest_0(isu_io_wb_rfDest_0),
    .io_wb_rfDest_1(isu_io_wb_rfDest_1),
    .io_wb_rfDest_2(isu_io_wb_rfDest_2),
    .io_wb_rfDest_3(isu_io_wb_rfDest_3),
    .io_wb_rfDest_4(isu_io_wb_rfDest_4),
    .io_wb_rfDest_5(isu_io_wb_rfDest_5),
    .io_wb_rfDest_6(isu_io_wb_rfDest_6),
    .io_wb_rfDest_7(isu_io_wb_rfDest_7),
    .io_wb_WriteData_0(isu_io_wb_WriteData_0),
    .io_wb_WriteData_1(isu_io_wb_WriteData_1),
    .io_wb_WriteData_2(isu_io_wb_WriteData_2),
    .io_wb_WriteData_3(isu_io_wb_WriteData_3),
    .io_wb_WriteData_4(isu_io_wb_WriteData_4),
    .io_wb_WriteData_5(isu_io_wb_WriteData_5),
    .io_wb_WriteData_6(isu_io_wb_WriteData_6),
    .io_wb_WriteData_7(isu_io_wb_WriteData_7),
    .io_wb_rfSrc1_0(isu_io_wb_rfSrc1_0),
    .io_wb_rfSrc1_1(isu_io_wb_rfSrc1_1),
    .io_wb_rfSrc2_0(isu_io_wb_rfSrc2_0),
    .io_wb_rfSrc2_1(isu_io_wb_rfSrc2_1),
    .io_wb_rfSrc3_0(isu_io_wb_rfSrc3_0),
    .io_wb_rfSrc3_1(isu_io_wb_rfSrc3_1),
    .io_wb_ReadData1_0(isu_io_wb_ReadData1_0),
    .io_wb_ReadData1_1(isu_io_wb_ReadData1_1),
    .io_wb_ReadData2_0(isu_io_wb_ReadData2_0),
    .io_wb_ReadData2_1(isu_io_wb_ReadData2_1),
    .io_wb_ReadData3_0(isu_io_wb_ReadData3_0),
    .io_wb_ReadData3_1(isu_io_wb_ReadData3_1),
    .io_wb_InstNo_0(isu_io_wb_InstNo_0),
    .io_wb_InstNo_1(isu_io_wb_InstNo_1),
    .io_wb_InstNo_2(isu_io_wb_InstNo_2),
    .io_wb_InstNo_3(isu_io_wb_InstNo_3),
    .io_wb_InstNo_4(isu_io_wb_InstNo_4),
    .io_wb_InstNo_5(isu_io_wb_InstNo_5),
    .io_wb_InstNo_6(isu_io_wb_InstNo_6),
    .io_wb_InstNo_7(isu_io_wb_InstNo_7),
    .io_forward_0_valid(isu_io_forward_0_valid),
    .io_forward_0_wb_rfWen(isu_io_forward_0_wb_rfWen),
    .io_forward_0_wb_rfDest(isu_io_forward_0_wb_rfDest),
    .io_forward_0_wb_rfData(isu_io_forward_0_wb_rfData),
    .io_forward_0_InstNo(isu_io_forward_0_InstNo),
    .io_forward_1_valid(isu_io_forward_1_valid),
    .io_forward_1_wb_rfWen(isu_io_forward_1_wb_rfWen),
    .io_forward_1_wb_rfDest(isu_io_forward_1_wb_rfDest),
    .io_forward_1_wb_rfData(isu_io_forward_1_wb_rfData),
    .io_forward_1_InstNo(isu_io_forward_1_InstNo),
    .io_forward_2_valid(isu_io_forward_2_valid),
    .io_forward_2_wb_rfWen(isu_io_forward_2_wb_rfWen),
    .io_forward_2_wb_rfDest(isu_io_forward_2_wb_rfDest),
    .io_forward_2_wb_rfData(isu_io_forward_2_wb_rfData),
    .io_forward_2_InstNo(isu_io_forward_2_InstNo),
    .io_forward_3_valid(isu_io_forward_3_valid),
    .io_forward_3_wb_rfWen(isu_io_forward_3_wb_rfWen),
    .io_forward_3_wb_rfDest(isu_io_forward_3_wb_rfDest),
    .io_forward_3_wb_rfData(isu_io_forward_3_wb_rfData),
    .io_forward_3_InstNo(isu_io_forward_3_InstNo),
    .io_forward_4_valid(isu_io_forward_4_valid),
    .io_forward_4_wb_rfWen(isu_io_forward_4_wb_rfWen),
    .io_forward_4_wb_rfDest(isu_io_forward_4_wb_rfDest),
    .io_forward_4_wb_rfData(isu_io_forward_4_wb_rfData),
    .io_forward_4_InstNo(isu_io_forward_4_InstNo),
    .io_forward_5_valid(isu_io_forward_5_valid),
    .io_forward_5_wb_rfWen(isu_io_forward_5_wb_rfWen),
    .io_forward_5_wb_rfDest(isu_io_forward_5_wb_rfDest),
    .io_forward_5_wb_rfData(isu_io_forward_5_wb_rfData),
    .io_forward_5_InstNo(isu_io_forward_5_InstNo),
    .io_forward_6_valid(isu_io_forward_6_valid),
    .io_forward_6_wb_rfWen(isu_io_forward_6_wb_rfWen),
    .io_forward_6_wb_rfDest(isu_io_forward_6_wb_rfDest),
    .io_forward_6_wb_rfData(isu_io_forward_6_wb_rfData),
    .io_forward_6_InstNo(isu_io_forward_6_InstNo),
    .io_forward_7_valid(isu_io_forward_7_valid),
    .io_forward_7_wb_rfWen(isu_io_forward_7_wb_rfWen),
    .io_forward_7_wb_rfDest(isu_io_forward_7_wb_rfDest),
    .io_forward_7_wb_rfData(isu_io_forward_7_wb_rfData),
    .io_forward_7_InstNo(isu_io_forward_7_InstNo),
    .io_flush(isu_io_flush),
    .io_num_enterwbu(isu_io_num_enterwbu),
    .io_TailPtr(isu_io_TailPtr)
  );
  new_SIMD_EXU exu ( // @[Backend.scala 725:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_0_ready(exu_io__in_0_ready),
    .io__in_0_valid(exu_io__in_0_valid),
    .io__in_0_bits_cf_instr(exu_io__in_0_bits_cf_instr),
    .io__in_0_bits_cf_pc(exu_io__in_0_bits_cf_pc),
    .io__in_0_bits_cf_pnpc(exu_io__in_0_bits_cf_pnpc),
    .io__in_0_bits_cf_brIdx(exu_io__in_0_bits_cf_brIdx),
    .io__in_0_bits_cf_runahead_checkpoint_id(exu_io__in_0_bits_cf_runahead_checkpoint_id),
    .io__in_0_bits_ctrl_fuOpType(exu_io__in_0_bits_ctrl_fuOpType),
    .io__in_0_bits_ctrl_rfWen(exu_io__in_0_bits_ctrl_rfWen),
    .io__in_0_bits_ctrl_rfDest(exu_io__in_0_bits_ctrl_rfDest),
    .io__in_0_bits_data_src1(exu_io__in_0_bits_data_src1),
    .io__in_0_bits_data_src2(exu_io__in_0_bits_data_src2),
    .io__in_0_bits_data_imm(exu_io__in_0_bits_data_imm),
    .io__in_0_bits_InstNo(exu_io__in_0_bits_InstNo),
    .io__in_0_bits_InstFlag(exu_io__in_0_bits_InstFlag),
    .io__in_1_ready(exu_io__in_1_ready),
    .io__in_1_valid(exu_io__in_1_valid),
    .io__in_1_bits_cf_pc(exu_io__in_1_bits_cf_pc),
    .io__in_1_bits_cf_exceptionVec_1(exu_io__in_1_bits_cf_exceptionVec_1),
    .io__in_1_bits_cf_exceptionVec_2(exu_io__in_1_bits_cf_exceptionVec_2),
    .io__in_1_bits_cf_exceptionVec_12(exu_io__in_1_bits_cf_exceptionVec_12),
    .io__in_1_bits_cf_intrVec_0(exu_io__in_1_bits_cf_intrVec_0),
    .io__in_1_bits_cf_intrVec_1(exu_io__in_1_bits_cf_intrVec_1),
    .io__in_1_bits_cf_intrVec_2(exu_io__in_1_bits_cf_intrVec_2),
    .io__in_1_bits_cf_intrVec_3(exu_io__in_1_bits_cf_intrVec_3),
    .io__in_1_bits_cf_intrVec_4(exu_io__in_1_bits_cf_intrVec_4),
    .io__in_1_bits_cf_intrVec_5(exu_io__in_1_bits_cf_intrVec_5),
    .io__in_1_bits_cf_intrVec_6(exu_io__in_1_bits_cf_intrVec_6),
    .io__in_1_bits_cf_intrVec_7(exu_io__in_1_bits_cf_intrVec_7),
    .io__in_1_bits_cf_intrVec_8(exu_io__in_1_bits_cf_intrVec_8),
    .io__in_1_bits_cf_intrVec_9(exu_io__in_1_bits_cf_intrVec_9),
    .io__in_1_bits_cf_intrVec_10(exu_io__in_1_bits_cf_intrVec_10),
    .io__in_1_bits_cf_intrVec_11(exu_io__in_1_bits_cf_intrVec_11),
    .io__in_1_bits_cf_crossPageIPFFix(exu_io__in_1_bits_cf_crossPageIPFFix),
    .io__in_1_bits_cf_runahead_checkpoint_id(exu_io__in_1_bits_cf_runahead_checkpoint_id),
    .io__in_1_bits_ctrl_fuOpType(exu_io__in_1_bits_ctrl_fuOpType),
    .io__in_1_bits_ctrl_rfWen(exu_io__in_1_bits_ctrl_rfWen),
    .io__in_1_bits_ctrl_rfDest(exu_io__in_1_bits_ctrl_rfDest),
    .io__in_1_bits_ctrl_isMou(exu_io__in_1_bits_ctrl_isMou),
    .io__in_1_bits_data_src1(exu_io__in_1_bits_data_src1),
    .io__in_1_bits_data_src2(exu_io__in_1_bits_data_src2),
    .io__in_1_bits_InstNo(exu_io__in_1_bits_InstNo),
    .io__in_1_bits_InstFlag(exu_io__in_1_bits_InstFlag),
    .io__in_2_ready(exu_io__in_2_ready),
    .io__in_2_valid(exu_io__in_2_valid),
    .io__in_2_bits_cf_instr(exu_io__in_2_bits_cf_instr),
    .io__in_2_bits_cf_pc(exu_io__in_2_bits_cf_pc),
    .io__in_2_bits_cf_runahead_checkpoint_id(exu_io__in_2_bits_cf_runahead_checkpoint_id),
    .io__in_2_bits_cf_instrType(exu_io__in_2_bits_cf_instrType),
    .io__in_2_bits_ctrl_fuOpType(exu_io__in_2_bits_ctrl_fuOpType),
    .io__in_2_bits_ctrl_funct3(exu_io__in_2_bits_ctrl_funct3),
    .io__in_2_bits_ctrl_func24(exu_io__in_2_bits_ctrl_func24),
    .io__in_2_bits_ctrl_func23(exu_io__in_2_bits_ctrl_func23),
    .io__in_2_bits_ctrl_rfWen(exu_io__in_2_bits_ctrl_rfWen),
    .io__in_2_bits_ctrl_rfDest(exu_io__in_2_bits_ctrl_rfDest),
    .io__in_2_bits_data_src1(exu_io__in_2_bits_data_src1),
    .io__in_2_bits_data_src2(exu_io__in_2_bits_data_src2),
    .io__in_2_bits_data_src3(exu_io__in_2_bits_data_src3),
    .io__in_2_bits_InstNo(exu_io__in_2_bits_InstNo),
    .io__in_2_bits_InstFlag(exu_io__in_2_bits_InstFlag),
    .io__in_3_ready(exu_io__in_3_ready),
    .io__in_3_valid(exu_io__in_3_valid),
    .io__in_3_bits_cf_instr(exu_io__in_3_bits_cf_instr),
    .io__in_3_bits_cf_pc(exu_io__in_3_bits_cf_pc),
    .io__in_3_bits_cf_runahead_checkpoint_id(exu_io__in_3_bits_cf_runahead_checkpoint_id),
    .io__in_3_bits_cf_instrType(exu_io__in_3_bits_cf_instrType),
    .io__in_3_bits_ctrl_fuOpType(exu_io__in_3_bits_ctrl_fuOpType),
    .io__in_3_bits_ctrl_funct3(exu_io__in_3_bits_ctrl_funct3),
    .io__in_3_bits_ctrl_func24(exu_io__in_3_bits_ctrl_func24),
    .io__in_3_bits_ctrl_func23(exu_io__in_3_bits_ctrl_func23),
    .io__in_3_bits_ctrl_rfWen(exu_io__in_3_bits_ctrl_rfWen),
    .io__in_3_bits_ctrl_rfDest(exu_io__in_3_bits_ctrl_rfDest),
    .io__in_3_bits_data_src1(exu_io__in_3_bits_data_src1),
    .io__in_3_bits_data_src2(exu_io__in_3_bits_data_src2),
    .io__in_3_bits_data_src3(exu_io__in_3_bits_data_src3),
    .io__in_3_bits_InstNo(exu_io__in_3_bits_InstNo),
    .io__in_3_bits_InstFlag(exu_io__in_3_bits_InstFlag),
    .io__in_4_ready(exu_io__in_4_ready),
    .io__in_4_valid(exu_io__in_4_valid),
    .io__in_4_bits_cf_instr(exu_io__in_4_bits_cf_instr),
    .io__in_4_bits_cf_pc(exu_io__in_4_bits_cf_pc),
    .io__in_4_bits_cf_exceptionVec_1(exu_io__in_4_bits_cf_exceptionVec_1),
    .io__in_4_bits_cf_exceptionVec_2(exu_io__in_4_bits_cf_exceptionVec_2),
    .io__in_4_bits_cf_exceptionVec_12(exu_io__in_4_bits_cf_exceptionVec_12),
    .io__in_4_bits_cf_intrVec_0(exu_io__in_4_bits_cf_intrVec_0),
    .io__in_4_bits_cf_intrVec_1(exu_io__in_4_bits_cf_intrVec_1),
    .io__in_4_bits_cf_intrVec_2(exu_io__in_4_bits_cf_intrVec_2),
    .io__in_4_bits_cf_intrVec_3(exu_io__in_4_bits_cf_intrVec_3),
    .io__in_4_bits_cf_intrVec_4(exu_io__in_4_bits_cf_intrVec_4),
    .io__in_4_bits_cf_intrVec_5(exu_io__in_4_bits_cf_intrVec_5),
    .io__in_4_bits_cf_intrVec_6(exu_io__in_4_bits_cf_intrVec_6),
    .io__in_4_bits_cf_intrVec_7(exu_io__in_4_bits_cf_intrVec_7),
    .io__in_4_bits_cf_intrVec_8(exu_io__in_4_bits_cf_intrVec_8),
    .io__in_4_bits_cf_intrVec_9(exu_io__in_4_bits_cf_intrVec_9),
    .io__in_4_bits_cf_intrVec_10(exu_io__in_4_bits_cf_intrVec_10),
    .io__in_4_bits_cf_intrVec_11(exu_io__in_4_bits_cf_intrVec_11),
    .io__in_4_bits_cf_crossPageIPFFix(exu_io__in_4_bits_cf_crossPageIPFFix),
    .io__in_4_bits_cf_runahead_checkpoint_id(exu_io__in_4_bits_cf_runahead_checkpoint_id),
    .io__in_4_bits_ctrl_fuOpType(exu_io__in_4_bits_ctrl_fuOpType),
    .io__in_4_bits_ctrl_rfWen(exu_io__in_4_bits_ctrl_rfWen),
    .io__in_4_bits_ctrl_rfDest(exu_io__in_4_bits_ctrl_rfDest),
    .io__in_4_bits_ctrl_isMou(exu_io__in_4_bits_ctrl_isMou),
    .io__in_4_bits_data_src1(exu_io__in_4_bits_data_src1),
    .io__in_4_bits_data_src2(exu_io__in_4_bits_data_src2),
    .io__in_4_bits_data_imm(exu_io__in_4_bits_data_imm),
    .io__in_4_bits_InstNo(exu_io__in_4_bits_InstNo),
    .io__in_4_bits_InstFlag(exu_io__in_4_bits_InstFlag),
    .io__in_5_ready(exu_io__in_5_ready),
    .io__in_5_valid(exu_io__in_5_valid),
    .io__in_5_bits_cf_pc(exu_io__in_5_bits_cf_pc),
    .io__in_5_bits_cf_runahead_checkpoint_id(exu_io__in_5_bits_cf_runahead_checkpoint_id),
    .io__in_5_bits_ctrl_fuOpType(exu_io__in_5_bits_ctrl_fuOpType),
    .io__in_5_bits_ctrl_rfWen(exu_io__in_5_bits_ctrl_rfWen),
    .io__in_5_bits_ctrl_rfDest(exu_io__in_5_bits_ctrl_rfDest),
    .io__in_5_bits_data_src1(exu_io__in_5_bits_data_src1),
    .io__in_5_bits_data_src2(exu_io__in_5_bits_data_src2),
    .io__in_5_bits_InstNo(exu_io__in_5_bits_InstNo),
    .io__in_6_ready(exu_io__in_6_ready),
    .io__in_6_valid(exu_io__in_6_valid),
    .io__in_6_bits_cf_instr(exu_io__in_6_bits_cf_instr),
    .io__in_6_bits_cf_pc(exu_io__in_6_bits_cf_pc),
    .io__in_6_bits_cf_pnpc(exu_io__in_6_bits_cf_pnpc),
    .io__in_6_bits_cf_brIdx(exu_io__in_6_bits_cf_brIdx),
    .io__in_6_bits_cf_runahead_checkpoint_id(exu_io__in_6_bits_cf_runahead_checkpoint_id),
    .io__in_6_bits_ctrl_fuOpType(exu_io__in_6_bits_ctrl_fuOpType),
    .io__in_6_bits_ctrl_rfWen(exu_io__in_6_bits_ctrl_rfWen),
    .io__in_6_bits_ctrl_rfDest(exu_io__in_6_bits_ctrl_rfDest),
    .io__in_6_bits_data_src1(exu_io__in_6_bits_data_src1),
    .io__in_6_bits_data_src2(exu_io__in_6_bits_data_src2),
    .io__in_6_bits_data_imm(exu_io__in_6_bits_data_imm),
    .io__in_6_bits_InstNo(exu_io__in_6_bits_InstNo),
    .io__in_7_ready(exu_io__in_7_ready),
    .io__in_7_valid(exu_io__in_7_valid),
    .io__in_7_bits_cf_instr(exu_io__in_7_bits_cf_instr),
    .io__in_7_bits_cf_pc(exu_io__in_7_bits_cf_pc),
    .io__in_7_bits_cf_pnpc(exu_io__in_7_bits_cf_pnpc),
    .io__in_7_bits_cf_brIdx(exu_io__in_7_bits_cf_brIdx),
    .io__in_7_bits_cf_runahead_checkpoint_id(exu_io__in_7_bits_cf_runahead_checkpoint_id),
    .io__in_7_bits_ctrl_fuOpType(exu_io__in_7_bits_ctrl_fuOpType),
    .io__in_7_bits_ctrl_rfWen(exu_io__in_7_bits_ctrl_rfWen),
    .io__in_7_bits_ctrl_rfDest(exu_io__in_7_bits_ctrl_rfDest),
    .io__in_7_bits_data_src1(exu_io__in_7_bits_data_src1),
    .io__in_7_bits_data_src2(exu_io__in_7_bits_data_src2),
    .io__in_7_bits_data_imm(exu_io__in_7_bits_data_imm),
    .io__in_7_bits_InstNo(exu_io__in_7_bits_InstNo),
    .io__out_0_ready(exu_io__out_0_ready),
    .io__out_0_valid(exu_io__out_0_valid),
    .io__out_0_bits_decode_cf_pc(exu_io__out_0_bits_decode_cf_pc),
    .io__out_0_bits_decode_cf_redirect_target(exu_io__out_0_bits_decode_cf_redirect_target),
    .io__out_0_bits_decode_cf_redirect_valid(exu_io__out_0_bits_decode_cf_redirect_valid),
    .io__out_0_bits_decode_cf_runahead_checkpoint_id(exu_io__out_0_bits_decode_cf_runahead_checkpoint_id),
    .io__out_0_bits_decode_ctrl_rfWen(exu_io__out_0_bits_decode_ctrl_rfWen),
    .io__out_0_bits_decode_ctrl_rfDest(exu_io__out_0_bits_decode_ctrl_rfDest),
    .io__out_0_bits_decode_InstNo(exu_io__out_0_bits_decode_InstNo),
    .io__out_0_bits_decode_InstFlag(exu_io__out_0_bits_decode_InstFlag),
    .io__out_0_bits_commits(exu_io__out_0_bits_commits),
    .io__out_1_ready(exu_io__out_1_ready),
    .io__out_1_valid(exu_io__out_1_valid),
    .io__out_1_bits_decode_cf_pc(exu_io__out_1_bits_decode_cf_pc),
    .io__out_1_bits_decode_cf_redirect_target(exu_io__out_1_bits_decode_cf_redirect_target),
    .io__out_1_bits_decode_cf_redirect_valid(exu_io__out_1_bits_decode_cf_redirect_valid),
    .io__out_1_bits_decode_cf_runahead_checkpoint_id(exu_io__out_1_bits_decode_cf_runahead_checkpoint_id),
    .io__out_1_bits_decode_ctrl_rfWen(exu_io__out_1_bits_decode_ctrl_rfWen),
    .io__out_1_bits_decode_ctrl_rfDest(exu_io__out_1_bits_decode_ctrl_rfDest),
    .io__out_1_bits_decode_InstNo(exu_io__out_1_bits_decode_InstNo),
    .io__out_1_bits_decode_InstFlag(exu_io__out_1_bits_decode_InstFlag),
    .io__out_1_bits_commits(exu_io__out_1_bits_commits),
    .io__out_2_ready(exu_io__out_2_ready),
    .io__out_2_valid(exu_io__out_2_valid),
    .io__out_2_bits_decode_cf_pc(exu_io__out_2_bits_decode_cf_pc),
    .io__out_2_bits_decode_cf_runahead_checkpoint_id(exu_io__out_2_bits_decode_cf_runahead_checkpoint_id),
    .io__out_2_bits_decode_ctrl_rfWen(exu_io__out_2_bits_decode_ctrl_rfWen),
    .io__out_2_bits_decode_ctrl_rfDest(exu_io__out_2_bits_decode_ctrl_rfDest),
    .io__out_2_bits_decode_pext_OV(exu_io__out_2_bits_decode_pext_OV),
    .io__out_2_bits_decode_InstNo(exu_io__out_2_bits_decode_InstNo),
    .io__out_2_bits_commits(exu_io__out_2_bits_commits),
    .io__out_3_ready(exu_io__out_3_ready),
    .io__out_3_valid(exu_io__out_3_valid),
    .io__out_3_bits_decode_cf_pc(exu_io__out_3_bits_decode_cf_pc),
    .io__out_3_bits_decode_cf_runahead_checkpoint_id(exu_io__out_3_bits_decode_cf_runahead_checkpoint_id),
    .io__out_3_bits_decode_ctrl_rfWen(exu_io__out_3_bits_decode_ctrl_rfWen),
    .io__out_3_bits_decode_ctrl_rfDest(exu_io__out_3_bits_decode_ctrl_rfDest),
    .io__out_3_bits_decode_pext_OV(exu_io__out_3_bits_decode_pext_OV),
    .io__out_3_bits_decode_InstNo(exu_io__out_3_bits_decode_InstNo),
    .io__out_3_bits_commits(exu_io__out_3_bits_commits),
    .io__out_4_ready(exu_io__out_4_ready),
    .io__out_4_valid(exu_io__out_4_valid),
    .io__out_4_bits_decode_cf_pc(exu_io__out_4_bits_decode_cf_pc),
    .io__out_4_bits_decode_cf_runahead_checkpoint_id(exu_io__out_4_bits_decode_cf_runahead_checkpoint_id),
    .io__out_4_bits_decode_ctrl_rfWen(exu_io__out_4_bits_decode_ctrl_rfWen),
    .io__out_4_bits_decode_ctrl_rfDest(exu_io__out_4_bits_decode_ctrl_rfDest),
    .io__out_4_bits_decode_InstNo(exu_io__out_4_bits_decode_InstNo),
    .io__out_4_bits_commits(exu_io__out_4_bits_commits),
    .io__out_5_ready(exu_io__out_5_ready),
    .io__out_5_valid(exu_io__out_5_valid),
    .io__out_5_bits_decode_cf_pc(exu_io__out_5_bits_decode_cf_pc),
    .io__out_5_bits_decode_cf_runahead_checkpoint_id(exu_io__out_5_bits_decode_cf_runahead_checkpoint_id),
    .io__out_5_bits_decode_ctrl_rfWen(exu_io__out_5_bits_decode_ctrl_rfWen),
    .io__out_5_bits_decode_ctrl_rfDest(exu_io__out_5_bits_decode_ctrl_rfDest),
    .io__out_5_bits_decode_InstNo(exu_io__out_5_bits_decode_InstNo),
    .io__out_5_bits_commits(exu_io__out_5_bits_commits),
    .io__out_6_ready(exu_io__out_6_ready),
    .io__out_6_valid(exu_io__out_6_valid),
    .io__out_6_bits_decode_cf_pc(exu_io__out_6_bits_decode_cf_pc),
    .io__out_6_bits_decode_cf_redirect_target(exu_io__out_6_bits_decode_cf_redirect_target),
    .io__out_6_bits_decode_cf_redirect_valid(exu_io__out_6_bits_decode_cf_redirect_valid),
    .io__out_6_bits_decode_cf_runahead_checkpoint_id(exu_io__out_6_bits_decode_cf_runahead_checkpoint_id),
    .io__out_6_bits_decode_ctrl_rfWen(exu_io__out_6_bits_decode_ctrl_rfWen),
    .io__out_6_bits_decode_ctrl_rfDest(exu_io__out_6_bits_decode_ctrl_rfDest),
    .io__out_6_bits_decode_InstNo(exu_io__out_6_bits_decode_InstNo),
    .io__out_6_bits_commits(exu_io__out_6_bits_commits),
    .io__out_7_ready(exu_io__out_7_ready),
    .io__out_7_valid(exu_io__out_7_valid),
    .io__out_7_bits_decode_cf_pc(exu_io__out_7_bits_decode_cf_pc),
    .io__out_7_bits_decode_cf_redirect_target(exu_io__out_7_bits_decode_cf_redirect_target),
    .io__out_7_bits_decode_cf_redirect_valid(exu_io__out_7_bits_decode_cf_redirect_valid),
    .io__out_7_bits_decode_cf_runahead_checkpoint_id(exu_io__out_7_bits_decode_cf_runahead_checkpoint_id),
    .io__out_7_bits_decode_ctrl_rfWen(exu_io__out_7_bits_decode_ctrl_rfWen),
    .io__out_7_bits_decode_ctrl_rfDest(exu_io__out_7_bits_decode_ctrl_rfDest),
    .io__out_7_bits_decode_InstNo(exu_io__out_7_bits_decode_InstNo),
    .io__out_7_bits_commits(exu_io__out_7_bits_commits),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_0_valid(exu_io__forward_0_valid),
    .io__forward_0_wb_rfWen(exu_io__forward_0_wb_rfWen),
    .io__forward_0_wb_rfDest(exu_io__forward_0_wb_rfDest),
    .io__forward_0_wb_rfData(exu_io__forward_0_wb_rfData),
    .io__forward_0_InstNo(exu_io__forward_0_InstNo),
    .io__forward_1_valid(exu_io__forward_1_valid),
    .io__forward_1_wb_rfWen(exu_io__forward_1_wb_rfWen),
    .io__forward_1_wb_rfDest(exu_io__forward_1_wb_rfDest),
    .io__forward_1_wb_rfData(exu_io__forward_1_wb_rfData),
    .io__forward_1_InstNo(exu_io__forward_1_InstNo),
    .io__forward_2_valid(exu_io__forward_2_valid),
    .io__forward_2_wb_rfWen(exu_io__forward_2_wb_rfWen),
    .io__forward_2_wb_rfDest(exu_io__forward_2_wb_rfDest),
    .io__forward_2_wb_rfData(exu_io__forward_2_wb_rfData),
    .io__forward_2_InstNo(exu_io__forward_2_InstNo),
    .io__forward_3_valid(exu_io__forward_3_valid),
    .io__forward_3_wb_rfWen(exu_io__forward_3_wb_rfWen),
    .io__forward_3_wb_rfDest(exu_io__forward_3_wb_rfDest),
    .io__forward_3_wb_rfData(exu_io__forward_3_wb_rfData),
    .io__forward_3_InstNo(exu_io__forward_3_InstNo),
    .io__forward_4_valid(exu_io__forward_4_valid),
    .io__forward_4_wb_rfWen(exu_io__forward_4_wb_rfWen),
    .io__forward_4_wb_rfDest(exu_io__forward_4_wb_rfDest),
    .io__forward_4_wb_rfData(exu_io__forward_4_wb_rfData),
    .io__forward_4_InstNo(exu_io__forward_4_InstNo),
    .io__forward_5_valid(exu_io__forward_5_valid),
    .io__forward_5_wb_rfWen(exu_io__forward_5_wb_rfWen),
    .io__forward_5_wb_rfDest(exu_io__forward_5_wb_rfDest),
    .io__forward_5_wb_rfData(exu_io__forward_5_wb_rfData),
    .io__forward_5_InstNo(exu_io__forward_5_InstNo),
    .io__forward_6_valid(exu_io__forward_6_valid),
    .io__forward_6_wb_rfWen(exu_io__forward_6_wb_rfWen),
    .io__forward_6_wb_rfDest(exu_io__forward_6_wb_rfDest),
    .io__forward_6_wb_rfData(exu_io__forward_6_wb_rfData),
    .io__forward_6_InstNo(exu_io__forward_6_InstNo),
    .io__forward_7_valid(exu_io__forward_7_valid),
    .io__forward_7_wb_rfWen(exu_io__forward_7_wb_rfWen),
    .io__forward_7_wb_rfDest(exu_io__forward_7_wb_rfDest),
    .io__forward_7_wb_rfData(exu_io__forward_7_wb_rfData),
    .io__forward_7_InstNo(exu_io__forward_7_InstNo),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_addr(exu_io__memMMU_dmem_addr),
    .lsu_firststage_fire(exu_lsu_firststage_fire),
    ._T_408(exu__T_408),
    ._T_137_0(exu__T_137_0),
    .flushICache(exu_flushICache),
    ._T_140_0(exu__T_140_0),
    .perfCnts_2(exu_perfCnts_2),
    ._WIRE_2_0(exu__WIRE_2_0),
    .satp(exu_satp),
    .bpuUpdateReq_valid(exu_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(exu_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(exu_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(exu_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(exu_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(exu_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(exu_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(exu_bpuUpdateReq_isRVC),
    .io_in_0_valid(exu_io_in_0_valid),
    .ismmio(exu_ismmio),
    ._WIRE_2_1(exu__WIRE_2_1),
    .io_extra_mtip(exu_io_extra_mtip),
    .amoReq(exu_amoReq),
    ._T_136_0(exu__T_136_0),
    .io_extra_meip_0(exu_io_extra_meip_0),
    ._T_139_0(exu__T_139_0),
    .vmEnable(exu_vmEnable),
    .intrVec(exu_intrVec),
    ._T_407(exu__T_407),
    ._WIRE_1_0(exu__WIRE_1_0),
    .io_extra_msip(exu_io_extra_msip),
    ._T_138_0(exu__T_138_0),
    .flushTLB(exu_flushTLB),
    ._T_135_0(exu__T_135_0)
  );
  new_SIMD_WBU wbu ( // @[Backend.scala 726:20]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io__in_0_valid(wbu_io__in_0_valid),
    .io__in_0_bits_decode_cf_pc(wbu_io__in_0_bits_decode_cf_pc),
    .io__in_0_bits_decode_cf_redirect_target(wbu_io__in_0_bits_decode_cf_redirect_target),
    .io__in_0_bits_decode_cf_redirect_valid(wbu_io__in_0_bits_decode_cf_redirect_valid),
    .io__in_0_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_0_bits_decode_cf_runahead_checkpoint_id),
    .io__in_0_bits_decode_ctrl_rfWen(wbu_io__in_0_bits_decode_ctrl_rfWen),
    .io__in_0_bits_decode_ctrl_rfDest(wbu_io__in_0_bits_decode_ctrl_rfDest),
    .io__in_0_bits_decode_pext_OV(wbu_io__in_0_bits_decode_pext_OV),
    .io__in_0_bits_decode_InstNo(wbu_io__in_0_bits_decode_InstNo),
    .io__in_0_bits_commits(wbu_io__in_0_bits_commits),
    .io__in_1_valid(wbu_io__in_1_valid),
    .io__in_1_bits_decode_cf_pc(wbu_io__in_1_bits_decode_cf_pc),
    .io__in_1_bits_decode_cf_redirect_target(wbu_io__in_1_bits_decode_cf_redirect_target),
    .io__in_1_bits_decode_cf_redirect_valid(wbu_io__in_1_bits_decode_cf_redirect_valid),
    .io__in_1_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_1_bits_decode_cf_runahead_checkpoint_id),
    .io__in_1_bits_decode_ctrl_rfWen(wbu_io__in_1_bits_decode_ctrl_rfWen),
    .io__in_1_bits_decode_ctrl_rfDest(wbu_io__in_1_bits_decode_ctrl_rfDest),
    .io__in_1_bits_decode_pext_OV(wbu_io__in_1_bits_decode_pext_OV),
    .io__in_1_bits_decode_InstNo(wbu_io__in_1_bits_decode_InstNo),
    .io__in_1_bits_commits(wbu_io__in_1_bits_commits),
    .io__in_2_valid(wbu_io__in_2_valid),
    .io__in_2_bits_decode_cf_pc(wbu_io__in_2_bits_decode_cf_pc),
    .io__in_2_bits_decode_cf_redirect_target(wbu_io__in_2_bits_decode_cf_redirect_target),
    .io__in_2_bits_decode_cf_redirect_valid(wbu_io__in_2_bits_decode_cf_redirect_valid),
    .io__in_2_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_2_bits_decode_cf_runahead_checkpoint_id),
    .io__in_2_bits_decode_ctrl_rfWen(wbu_io__in_2_bits_decode_ctrl_rfWen),
    .io__in_2_bits_decode_ctrl_rfDest(wbu_io__in_2_bits_decode_ctrl_rfDest),
    .io__in_2_bits_decode_pext_OV(wbu_io__in_2_bits_decode_pext_OV),
    .io__in_2_bits_decode_InstNo(wbu_io__in_2_bits_decode_InstNo),
    .io__in_2_bits_commits(wbu_io__in_2_bits_commits),
    .io__in_3_valid(wbu_io__in_3_valid),
    .io__in_3_bits_decode_cf_pc(wbu_io__in_3_bits_decode_cf_pc),
    .io__in_3_bits_decode_cf_redirect_target(wbu_io__in_3_bits_decode_cf_redirect_target),
    .io__in_3_bits_decode_cf_redirect_valid(wbu_io__in_3_bits_decode_cf_redirect_valid),
    .io__in_3_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_3_bits_decode_cf_runahead_checkpoint_id),
    .io__in_3_bits_decode_ctrl_rfWen(wbu_io__in_3_bits_decode_ctrl_rfWen),
    .io__in_3_bits_decode_ctrl_rfDest(wbu_io__in_3_bits_decode_ctrl_rfDest),
    .io__in_3_bits_decode_pext_OV(wbu_io__in_3_bits_decode_pext_OV),
    .io__in_3_bits_decode_InstNo(wbu_io__in_3_bits_decode_InstNo),
    .io__in_3_bits_commits(wbu_io__in_3_bits_commits),
    .io__in_4_valid(wbu_io__in_4_valid),
    .io__in_4_bits_decode_cf_pc(wbu_io__in_4_bits_decode_cf_pc),
    .io__in_4_bits_decode_cf_redirect_target(wbu_io__in_4_bits_decode_cf_redirect_target),
    .io__in_4_bits_decode_cf_redirect_valid(wbu_io__in_4_bits_decode_cf_redirect_valid),
    .io__in_4_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_4_bits_decode_cf_runahead_checkpoint_id),
    .io__in_4_bits_decode_ctrl_rfWen(wbu_io__in_4_bits_decode_ctrl_rfWen),
    .io__in_4_bits_decode_ctrl_rfDest(wbu_io__in_4_bits_decode_ctrl_rfDest),
    .io__in_4_bits_decode_pext_OV(wbu_io__in_4_bits_decode_pext_OV),
    .io__in_4_bits_decode_InstNo(wbu_io__in_4_bits_decode_InstNo),
    .io__in_4_bits_commits(wbu_io__in_4_bits_commits),
    .io__in_5_valid(wbu_io__in_5_valid),
    .io__in_5_bits_decode_cf_pc(wbu_io__in_5_bits_decode_cf_pc),
    .io__in_5_bits_decode_cf_redirect_target(wbu_io__in_5_bits_decode_cf_redirect_target),
    .io__in_5_bits_decode_cf_redirect_valid(wbu_io__in_5_bits_decode_cf_redirect_valid),
    .io__in_5_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_5_bits_decode_cf_runahead_checkpoint_id),
    .io__in_5_bits_decode_ctrl_rfWen(wbu_io__in_5_bits_decode_ctrl_rfWen),
    .io__in_5_bits_decode_ctrl_rfDest(wbu_io__in_5_bits_decode_ctrl_rfDest),
    .io__in_5_bits_decode_pext_OV(wbu_io__in_5_bits_decode_pext_OV),
    .io__in_5_bits_decode_InstNo(wbu_io__in_5_bits_decode_InstNo),
    .io__in_5_bits_commits(wbu_io__in_5_bits_commits),
    .io__in_6_valid(wbu_io__in_6_valid),
    .io__in_6_bits_decode_cf_pc(wbu_io__in_6_bits_decode_cf_pc),
    .io__in_6_bits_decode_cf_redirect_target(wbu_io__in_6_bits_decode_cf_redirect_target),
    .io__in_6_bits_decode_cf_redirect_valid(wbu_io__in_6_bits_decode_cf_redirect_valid),
    .io__in_6_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_6_bits_decode_cf_runahead_checkpoint_id),
    .io__in_6_bits_decode_ctrl_rfWen(wbu_io__in_6_bits_decode_ctrl_rfWen),
    .io__in_6_bits_decode_ctrl_rfDest(wbu_io__in_6_bits_decode_ctrl_rfDest),
    .io__in_6_bits_decode_pext_OV(wbu_io__in_6_bits_decode_pext_OV),
    .io__in_6_bits_decode_InstNo(wbu_io__in_6_bits_decode_InstNo),
    .io__in_6_bits_commits(wbu_io__in_6_bits_commits),
    .io__in_7_valid(wbu_io__in_7_valid),
    .io__in_7_bits_decode_cf_pc(wbu_io__in_7_bits_decode_cf_pc),
    .io__in_7_bits_decode_cf_redirect_target(wbu_io__in_7_bits_decode_cf_redirect_target),
    .io__in_7_bits_decode_cf_redirect_valid(wbu_io__in_7_bits_decode_cf_redirect_valid),
    .io__in_7_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_7_bits_decode_cf_runahead_checkpoint_id),
    .io__in_7_bits_decode_ctrl_rfWen(wbu_io__in_7_bits_decode_ctrl_rfWen),
    .io__in_7_bits_decode_ctrl_rfDest(wbu_io__in_7_bits_decode_ctrl_rfDest),
    .io__in_7_bits_decode_pext_OV(wbu_io__in_7_bits_decode_pext_OV),
    .io__in_7_bits_decode_InstNo(wbu_io__in_7_bits_decode_InstNo),
    .io__in_7_bits_commits(wbu_io__in_7_bits_commits),
    .io__wb_rfWen_0(wbu_io__wb_rfWen_0),
    .io__wb_rfWen_1(wbu_io__wb_rfWen_1),
    .io__wb_rfWen_2(wbu_io__wb_rfWen_2),
    .io__wb_rfWen_3(wbu_io__wb_rfWen_3),
    .io__wb_rfWen_4(wbu_io__wb_rfWen_4),
    .io__wb_rfWen_5(wbu_io__wb_rfWen_5),
    .io__wb_rfWen_6(wbu_io__wb_rfWen_6),
    .io__wb_rfWen_7(wbu_io__wb_rfWen_7),
    .io__wb_rfDest_0(wbu_io__wb_rfDest_0),
    .io__wb_rfDest_1(wbu_io__wb_rfDest_1),
    .io__wb_rfDest_2(wbu_io__wb_rfDest_2),
    .io__wb_rfDest_3(wbu_io__wb_rfDest_3),
    .io__wb_rfDest_4(wbu_io__wb_rfDest_4),
    .io__wb_rfDest_5(wbu_io__wb_rfDest_5),
    .io__wb_rfDest_6(wbu_io__wb_rfDest_6),
    .io__wb_rfDest_7(wbu_io__wb_rfDest_7),
    .io__wb_WriteData_0(wbu_io__wb_WriteData_0),
    .io__wb_WriteData_1(wbu_io__wb_WriteData_1),
    .io__wb_WriteData_2(wbu_io__wb_WriteData_2),
    .io__wb_WriteData_3(wbu_io__wb_WriteData_3),
    .io__wb_WriteData_4(wbu_io__wb_WriteData_4),
    .io__wb_WriteData_5(wbu_io__wb_WriteData_5),
    .io__wb_WriteData_6(wbu_io__wb_WriteData_6),
    .io__wb_WriteData_7(wbu_io__wb_WriteData_7),
    .io__wb_rfSrc1_0(wbu_io__wb_rfSrc1_0),
    .io__wb_rfSrc1_1(wbu_io__wb_rfSrc1_1),
    .io__wb_rfSrc2_0(wbu_io__wb_rfSrc2_0),
    .io__wb_rfSrc2_1(wbu_io__wb_rfSrc2_1),
    .io__wb_rfSrc3_0(wbu_io__wb_rfSrc3_0),
    .io__wb_rfSrc3_1(wbu_io__wb_rfSrc3_1),
    .io__wb_ReadData1_0(wbu_io__wb_ReadData1_0),
    .io__wb_ReadData1_1(wbu_io__wb_ReadData1_1),
    .io__wb_ReadData2_0(wbu_io__wb_ReadData2_0),
    .io__wb_ReadData2_1(wbu_io__wb_ReadData2_1),
    .io__wb_ReadData3_0(wbu_io__wb_ReadData3_0),
    .io__wb_ReadData3_1(wbu_io__wb_ReadData3_1),
    .io__wb_InstNo_0(wbu_io__wb_InstNo_0),
    .io__wb_InstNo_1(wbu_io__wb_InstNo_1),
    .io__wb_InstNo_2(wbu_io__wb_InstNo_2),
    .io__wb_InstNo_3(wbu_io__wb_InstNo_3),
    .io__wb_InstNo_4(wbu_io__wb_InstNo_4),
    .io__wb_InstNo_5(wbu_io__wb_InstNo_5),
    .io__wb_InstNo_6(wbu_io__wb_InstNo_6),
    .io__wb_InstNo_7(wbu_io__wb_InstNo_7),
    .io__redirect_valid(wbu_io__redirect_valid),
    ._T_137_0(wbu__T_137_0),
    ._T_140_0(wbu__T_140_0),
    .io_in_0_bits_decode_cf_pc(wbu_io_in_0_bits_decode_cf_pc),
    .io_wb_rfDest_0(wbu_io_wb_rfDest_0),
    .io_in_0_valid(wbu_io_in_0_valid),
    ._WIRE_2_1(wbu__WIRE_2_1),
    ._T_136_0(wbu__T_136_0),
    ._T_139_0(wbu__T_139_0),
    .io_wb_rfWen_0(wbu_io_wb_rfWen_0),
    .io_wb_WriteData_0(wbu_io_wb_WriteData_0),
    ._T_138_0(wbu__T_138_0),
    .io_in_0_valid_0(wbu_io_in_0_valid_0),
    ._T_135_0(wbu__T_135_0)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[Backend.scala 892:13]
  assign io_in_1_ready = isu_io_in_1_ready; // @[Backend.scala 892:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[Backend.scala 933:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[Backend.scala 933:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[Backend.scala 933:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[Backend.scala 933:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[Backend.scala 933:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[Backend.scala 933:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 931:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 932:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[Backend.scala 932:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 932:18]
  assign io_redirect_target = 3'h7 == _GEN_5930 ? exu_io__out_7_bits_decode_cf_redirect_target : _GEN_5774; // @[]
  assign io_redirect_valid = _GEN_5759 & _T_2274; // @[Backend.scala 924:77]
  assign flushICache = exu_flushICache;
  assign perfCnts_2 = exu_perfCnts_2;
  assign io_in_0_bits_decode_cf_pc = wbu_io_in_0_bits_decode_cf_pc;
  assign satp = exu_satp;
  assign bpuUpdateReq_valid = exu_bpuUpdateReq_valid;
  assign bpuUpdateReq_pc = exu_bpuUpdateReq_pc;
  assign bpuUpdateReq_isMissPredict = exu_bpuUpdateReq_isMissPredict;
  assign bpuUpdateReq_actualTarget = exu_bpuUpdateReq_actualTarget;
  assign bpuUpdateReq_actualTaken = exu_bpuUpdateReq_actualTaken;
  assign bpuUpdateReq_fuOpType = exu_bpuUpdateReq_fuOpType;
  assign bpuUpdateReq_btbType = exu_bpuUpdateReq_btbType;
  assign bpuUpdateReq_isRVC = exu_bpuUpdateReq_isRVC;
  assign io_wb_rfDest_0 = wbu_io_wb_rfDest_0;
  assign amoReq = exu_amoReq;
  assign io_wb_rfWen_0 = wbu_io_wb_rfWen_0;
  assign io_wb_WriteData_0 = wbu_io_wb_WriteData_0;
  assign intrVec = exu_intrVec;
  assign flushTLB = exu_flushTLB;
  assign io_in_0_valid_0 = wbu_io_in_0_valid_0;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_runahead_checkpoint_id = io_in_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_cf_instrType = io_in_0_bits_cf_instrType; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_funct3 = io_in_0_bits_ctrl_funct3; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_func24 = io_in_0_bits_ctrl_func24; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_func23 = io_in_0_bits_ctrl_func23; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_rfSrc3 = io_in_0_bits_ctrl_rfSrc3; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_ctrl_isMou = io_in_0_bits_ctrl_isMou; // @[Backend.scala 892:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[Backend.scala 892:13]
  assign isu_io_in_1_valid = io_in_1_valid; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_instr = io_in_1_bits_cf_instr; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_pc = io_in_1_bits_cf_pc; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_pnpc = io_in_1_bits_cf_pnpc; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_exceptionVec_1 = io_in_1_bits_cf_exceptionVec_1; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_exceptionVec_2 = io_in_1_bits_cf_exceptionVec_2; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_exceptionVec_12 = io_in_1_bits_cf_exceptionVec_12; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_0 = io_in_1_bits_cf_intrVec_0; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_1 = io_in_1_bits_cf_intrVec_1; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_2 = io_in_1_bits_cf_intrVec_2; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_3 = io_in_1_bits_cf_intrVec_3; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_4 = io_in_1_bits_cf_intrVec_4; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_5 = io_in_1_bits_cf_intrVec_5; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_6 = io_in_1_bits_cf_intrVec_6; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_7 = io_in_1_bits_cf_intrVec_7; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_8 = io_in_1_bits_cf_intrVec_8; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_9 = io_in_1_bits_cf_intrVec_9; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_10 = io_in_1_bits_cf_intrVec_10; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_intrVec_11 = io_in_1_bits_cf_intrVec_11; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_brIdx = io_in_1_bits_cf_brIdx; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_crossPageIPFFix = io_in_1_bits_cf_crossPageIPFFix; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_runahead_checkpoint_id = io_in_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_cf_instrType = io_in_1_bits_cf_instrType; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_src1Type = io_in_1_bits_ctrl_src1Type; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_src2Type = io_in_1_bits_ctrl_src2Type; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_fuType = io_in_1_bits_ctrl_fuType; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_fuOpType = io_in_1_bits_ctrl_fuOpType; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_funct3 = io_in_1_bits_ctrl_funct3; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_func24 = io_in_1_bits_ctrl_func24; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_func23 = io_in_1_bits_ctrl_func23; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_rfSrc1 = io_in_1_bits_ctrl_rfSrc1; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_rfSrc2 = io_in_1_bits_ctrl_rfSrc2; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_rfSrc3 = io_in_1_bits_ctrl_rfSrc3; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_rfWen = io_in_1_bits_ctrl_rfWen; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_rfDest = io_in_1_bits_ctrl_rfDest; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_ctrl_isMou = io_in_1_bits_ctrl_isMou; // @[Backend.scala 892:13]
  assign isu_io_in_1_bits_data_imm = io_in_1_bits_data_imm; // @[Backend.scala 892:13]
  assign isu_io_out_0_ready = match_operaotr_0_7 | (match_operaotr_0_6 | (match_operaotr_0_5 | (match_operaotr_0_4 | (
    match_operaotr_0_3 | (match_operaotr_0_2 | (match_operaotr_0_1 | match_operaotr_0_0)))))); // @[Backend.scala 805:244 807:31]
  assign isu_io_out_1_ready = match_operaotr_1_7 | (match_operaotr_1_6 | (match_operaotr_1_5 | (match_operaotr_1_4 | (
    match_operaotr_1_3 | (match_operaotr_1_2 | (match_operaotr_1_1 | match_operaotr_1_0)))))); // @[Backend.scala 805:244 807:31]
  assign isu_io_wb_rfWen_0 = wbu_io__wb_rfWen_0; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_1 = wbu_io__wb_rfWen_1; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_2 = wbu_io__wb_rfWen_2; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_3 = wbu_io__wb_rfWen_3; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_4 = wbu_io__wb_rfWen_4; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_5 = wbu_io__wb_rfWen_5; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_6 = wbu_io__wb_rfWen_6; // @[Backend.scala 905:24]
  assign isu_io_wb_rfWen_7 = wbu_io__wb_rfWen_7; // @[Backend.scala 905:24]
  assign isu_io_wb_rfDest_0 = wbu_io__wb_rfDest_0; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_1 = wbu_io__wb_rfDest_1; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_2 = wbu_io__wb_rfDest_2; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_3 = wbu_io__wb_rfDest_3; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_4 = wbu_io__wb_rfDest_4; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_5 = wbu_io__wb_rfDest_5; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_6 = wbu_io__wb_rfDest_6; // @[Backend.scala 906:24]
  assign isu_io_wb_rfDest_7 = wbu_io__wb_rfDest_7; // @[Backend.scala 906:24]
  assign isu_io_wb_WriteData_0 = wbu_io__wb_WriteData_0; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_1 = wbu_io__wb_WriteData_1; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_2 = wbu_io__wb_WriteData_2; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_3 = wbu_io__wb_WriteData_3; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_4 = wbu_io__wb_WriteData_4; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_5 = wbu_io__wb_WriteData_5; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_6 = wbu_io__wb_WriteData_6; // @[Backend.scala 907:27]
  assign isu_io_wb_WriteData_7 = wbu_io__wb_WriteData_7; // @[Backend.scala 907:27]
  assign isu_io_wb_ReadData1_0 = wbu_io__wb_ReadData1_0; // @[Backend.scala 912:27]
  assign isu_io_wb_ReadData1_1 = wbu_io__wb_ReadData1_1; // @[Backend.scala 912:27]
  assign isu_io_wb_ReadData2_0 = wbu_io__wb_ReadData2_0; // @[Backend.scala 913:27]
  assign isu_io_wb_ReadData2_1 = wbu_io__wb_ReadData2_1; // @[Backend.scala 913:27]
  assign isu_io_wb_ReadData3_0 = wbu_io__wb_ReadData3_0; // @[Backend.scala 919:29]
  assign isu_io_wb_ReadData3_1 = wbu_io__wb_ReadData3_1; // @[Backend.scala 919:29]
  assign isu_io_wb_InstNo_0 = wbu_io__wb_InstNo_0; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_1 = wbu_io__wb_InstNo_1; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_2 = wbu_io__wb_InstNo_2; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_3 = wbu_io__wb_InstNo_3; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_4 = wbu_io__wb_InstNo_4; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_5 = wbu_io__wb_InstNo_5; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_6 = wbu_io__wb_InstNo_6; // @[Backend.scala 909:24]
  assign isu_io_wb_InstNo_7 = wbu_io__wb_InstNo_7; // @[Backend.scala 909:24]
  assign isu_io_forward_0_valid = exu_io__forward_0_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_0_wb_rfWen = exu_io__forward_0_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_0_wb_rfDest = exu_io__forward_0_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_0_wb_rfData = exu_io__forward_0_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_0_InstNo = exu_io__forward_0_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_1_valid = exu_io__forward_1_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_1_wb_rfWen = exu_io__forward_1_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_1_wb_rfDest = exu_io__forward_1_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_1_wb_rfData = exu_io__forward_1_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_1_InstNo = exu_io__forward_1_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_2_valid = exu_io__forward_2_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_2_wb_rfWen = exu_io__forward_2_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_2_wb_rfDest = exu_io__forward_2_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_2_wb_rfData = exu_io__forward_2_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_2_InstNo = exu_io__forward_2_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_3_valid = exu_io__forward_3_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_3_wb_rfWen = exu_io__forward_3_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_3_wb_rfDest = exu_io__forward_3_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_3_wb_rfData = exu_io__forward_3_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_3_InstNo = exu_io__forward_3_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_4_valid = exu_io__forward_4_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_4_wb_rfWen = exu_io__forward_4_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_4_wb_rfDest = exu_io__forward_4_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_4_wb_rfData = exu_io__forward_4_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_4_InstNo = exu_io__forward_4_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_5_valid = exu_io__forward_5_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_5_wb_rfWen = exu_io__forward_5_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_5_wb_rfDest = exu_io__forward_5_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_5_wb_rfData = exu_io__forward_5_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_5_InstNo = exu_io__forward_5_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_6_valid = exu_io__forward_6_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_6_wb_rfWen = exu_io__forward_6_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_6_wb_rfDest = exu_io__forward_6_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_6_wb_rfData = exu_io__forward_6_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_6_InstNo = exu_io__forward_6_InstNo; // @[Backend.scala 928:23]
  assign isu_io_forward_7_valid = exu_io__forward_7_valid; // @[Backend.scala 928:23]
  assign isu_io_forward_7_wb_rfWen = exu_io__forward_7_wb_rfWen; // @[Backend.scala 928:23]
  assign isu_io_forward_7_wb_rfDest = exu_io__forward_7_wb_rfDest; // @[Backend.scala 928:23]
  assign isu_io_forward_7_wb_rfData = exu_io__forward_7_wb_rfData; // @[Backend.scala 928:23]
  assign isu_io_forward_7_InstNo = exu_io__forward_7_InstNo; // @[Backend.scala 928:23]
  assign isu_io_flush = io_flush[0]; // @[Backend.scala 901:27]
  assign isu_io_num_enterwbu = num_enterwbu[4:0]; // @[Backend.scala 899:23]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_0_valid = exu_valid_0; // @[Backend.scala 771:24]
  assign exu_io__in_0_bits_cf_instr = exu_bits_0_cf_instr; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_cf_pc = exu_bits_0_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_cf_pnpc = exu_bits_0_cf_pnpc; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_cf_brIdx = exu_bits_0_cf_brIdx; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_cf_runahead_checkpoint_id = exu_bits_0_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_ctrl_fuOpType = exu_bits_0_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_ctrl_rfWen = exu_bits_0_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_ctrl_rfDest = exu_bits_0_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_data_src1 = exu_bits_0_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_data_src2 = exu_bits_0_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_data_imm = exu_bits_0_data_imm; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_InstNo = exu_bits_0_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_0_bits_InstFlag = exu_bits_0_InstFlag; // @[Backend.scala 770:23]
  assign exu_io__in_1_valid = exu_valid_1; // @[Backend.scala 771:24]
  assign exu_io__in_1_bits_cf_pc = exu_bits_1_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_exceptionVec_1 = exu_bits_1_cf_exceptionVec_1; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_exceptionVec_2 = exu_bits_1_cf_exceptionVec_2; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_exceptionVec_12 = exu_bits_1_cf_exceptionVec_12; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_0 = exu_bits_1_cf_intrVec_0; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_1 = exu_bits_1_cf_intrVec_1; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_2 = exu_bits_1_cf_intrVec_2; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_3 = exu_bits_1_cf_intrVec_3; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_4 = exu_bits_1_cf_intrVec_4; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_5 = exu_bits_1_cf_intrVec_5; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_6 = exu_bits_1_cf_intrVec_6; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_7 = exu_bits_1_cf_intrVec_7; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_8 = exu_bits_1_cf_intrVec_8; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_9 = exu_bits_1_cf_intrVec_9; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_10 = exu_bits_1_cf_intrVec_10; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_intrVec_11 = exu_bits_1_cf_intrVec_11; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_crossPageIPFFix = exu_bits_1_cf_crossPageIPFFix; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_cf_runahead_checkpoint_id = exu_bits_1_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_ctrl_fuOpType = exu_bits_1_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_ctrl_rfWen = exu_bits_1_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_ctrl_rfDest = exu_bits_1_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_ctrl_isMou = exu_bits_1_ctrl_isMou; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_data_src1 = exu_bits_1_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_data_src2 = exu_bits_1_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_InstNo = exu_bits_1_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_1_bits_InstFlag = exu_bits_1_InstFlag; // @[Backend.scala 770:23]
  assign exu_io__in_2_valid = exu_valid_2; // @[Backend.scala 771:24]
  assign exu_io__in_2_bits_cf_instr = exu_bits_2_cf_instr; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_cf_pc = exu_bits_2_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_cf_runahead_checkpoint_id = exu_bits_2_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_cf_instrType = exu_bits_2_cf_instrType; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_ctrl_fuOpType = exu_bits_2_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_ctrl_funct3 = exu_bits_2_ctrl_funct3; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_ctrl_func24 = exu_bits_2_ctrl_func24; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_ctrl_func23 = exu_bits_2_ctrl_func23; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_ctrl_rfWen = exu_bits_2_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_ctrl_rfDest = exu_bits_2_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_data_src1 = exu_bits_2_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_data_src2 = exu_bits_2_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_data_src3 = exu_bits_2_data_src3; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_InstNo = exu_bits_2_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_2_bits_InstFlag = exu_bits_2_InstFlag; // @[Backend.scala 770:23]
  assign exu_io__in_3_valid = exu_valid_3; // @[Backend.scala 771:24]
  assign exu_io__in_3_bits_cf_instr = exu_bits_3_cf_instr; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_cf_pc = exu_bits_3_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_cf_runahead_checkpoint_id = exu_bits_3_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_cf_instrType = exu_bits_3_cf_instrType; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_ctrl_fuOpType = exu_bits_3_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_ctrl_funct3 = exu_bits_3_ctrl_funct3; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_ctrl_func24 = exu_bits_3_ctrl_func24; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_ctrl_func23 = exu_bits_3_ctrl_func23; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_ctrl_rfWen = exu_bits_3_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_ctrl_rfDest = exu_bits_3_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_data_src1 = exu_bits_3_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_data_src2 = exu_bits_3_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_data_src3 = exu_bits_3_data_src3; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_InstNo = exu_bits_3_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_3_bits_InstFlag = exu_bits_3_InstFlag; // @[Backend.scala 770:23]
  assign exu_io__in_4_valid = exu_valid_4; // @[Backend.scala 771:24]
  assign exu_io__in_4_bits_cf_instr = exu_bits_4_cf_instr; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_pc = exu_bits_4_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_exceptionVec_1 = exu_bits_4_cf_exceptionVec_1; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_exceptionVec_2 = exu_bits_4_cf_exceptionVec_2; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_exceptionVec_12 = exu_bits_4_cf_exceptionVec_12; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_0 = exu_bits_4_cf_intrVec_0; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_1 = exu_bits_4_cf_intrVec_1; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_2 = exu_bits_4_cf_intrVec_2; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_3 = exu_bits_4_cf_intrVec_3; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_4 = exu_bits_4_cf_intrVec_4; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_5 = exu_bits_4_cf_intrVec_5; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_6 = exu_bits_4_cf_intrVec_6; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_7 = exu_bits_4_cf_intrVec_7; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_8 = exu_bits_4_cf_intrVec_8; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_9 = exu_bits_4_cf_intrVec_9; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_10 = exu_bits_4_cf_intrVec_10; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_intrVec_11 = exu_bits_4_cf_intrVec_11; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_crossPageIPFFix = exu_bits_4_cf_crossPageIPFFix; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_cf_runahead_checkpoint_id = exu_bits_4_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_ctrl_fuOpType = exu_bits_4_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_ctrl_rfWen = exu_bits_4_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_ctrl_rfDest = exu_bits_4_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_ctrl_isMou = exu_bits_4_ctrl_isMou; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_data_src1 = exu_bits_4_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_data_src2 = exu_bits_4_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_data_imm = exu_bits_4_data_imm; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_InstNo = exu_bits_4_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_4_bits_InstFlag = exu_bits_4_InstFlag; // @[Backend.scala 770:23]
  assign exu_io__in_5_valid = exu_valid_5; // @[Backend.scala 771:24]
  assign exu_io__in_5_bits_cf_pc = exu_bits_5_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_cf_runahead_checkpoint_id = exu_bits_5_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_ctrl_fuOpType = exu_bits_5_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_ctrl_rfWen = exu_bits_5_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_ctrl_rfDest = exu_bits_5_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_data_src1 = exu_bits_5_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_data_src2 = exu_bits_5_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_5_bits_InstNo = exu_bits_5_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_6_valid = exu_valid_6; // @[Backend.scala 771:24]
  assign exu_io__in_6_bits_cf_instr = exu_bits_6_cf_instr; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_cf_pc = exu_bits_6_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_cf_pnpc = exu_bits_6_cf_pnpc; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_cf_brIdx = exu_bits_6_cf_brIdx; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_cf_runahead_checkpoint_id = exu_bits_6_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_ctrl_fuOpType = exu_bits_6_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_ctrl_rfWen = exu_bits_6_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_ctrl_rfDest = exu_bits_6_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_data_src1 = exu_bits_6_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_data_src2 = exu_bits_6_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_data_imm = exu_bits_6_data_imm; // @[Backend.scala 770:23]
  assign exu_io__in_6_bits_InstNo = exu_bits_6_InstNo; // @[Backend.scala 770:23]
  assign exu_io__in_7_valid = exu_valid_7; // @[Backend.scala 771:24]
  assign exu_io__in_7_bits_cf_instr = exu_bits_7_cf_instr; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_cf_pc = exu_bits_7_cf_pc; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_cf_pnpc = exu_bits_7_cf_pnpc; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_cf_brIdx = exu_bits_7_cf_brIdx; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_cf_runahead_checkpoint_id = exu_bits_7_cf_runahead_checkpoint_id; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_ctrl_fuOpType = exu_bits_7_ctrl_fuOpType; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_ctrl_rfWen = exu_bits_7_ctrl_rfWen; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_ctrl_rfDest = exu_bits_7_ctrl_rfDest; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_data_src1 = exu_bits_7_data_src1; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_data_src2 = exu_bits_7_data_src2; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_data_imm = exu_bits_7_data_imm; // @[Backend.scala 770:23]
  assign exu_io__in_7_bits_InstNo = exu_bits_7_InstNo; // @[Backend.scala 770:23]
  assign exu_io__out_0_ready = match_exuwbu_7_0 | (match_exuwbu_6_0 | (match_exuwbu_5_0 | (match_exuwbu_4_0 | (
    match_exuwbu_3_0 | (match_exuwbu_2_0 | (match_exuwbu_1_0 | match_exuwbu_0_0)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__out_1_ready = match_exuwbu_7_1 | (match_exuwbu_6_1 | (match_exuwbu_5_1 | (match_exuwbu_4_1 | (
    match_exuwbu_3_1 | (match_exuwbu_2_1 | (match_exuwbu_1_1 | match_exuwbu_0_1)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__out_2_ready = match_exuwbu_7_2 | (match_exuwbu_6_2 | (match_exuwbu_5_2 | (match_exuwbu_4_2 | (
    match_exuwbu_3_2 | (match_exuwbu_2_2 | (match_exuwbu_1_2 | match_exuwbu_0_2)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__out_3_ready = match_exuwbu_7_3 | (match_exuwbu_6_3 | (match_exuwbu_5_3 | (match_exuwbu_4_3 | (
    match_exuwbu_3_3 | (match_exuwbu_2_3 | (match_exuwbu_1_3 | match_exuwbu_0_3)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__out_4_ready = 6'h7 < lsuInstNo & ~wbu_valid_next_7 ? 1'h0 : _GEN_5742; // @[Backend.scala 878:48 879:19]
  assign exu_io__out_5_ready = match_exuwbu_7_5 | (match_exuwbu_6_5 | (match_exuwbu_5_5 | (match_exuwbu_4_5 | (
    match_exuwbu_3_5 | (match_exuwbu_2_5 | (match_exuwbu_1_5 | match_exuwbu_0_5)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__out_6_ready = match_exuwbu_7_6 | (match_exuwbu_6_6 | (match_exuwbu_5_6 | (match_exuwbu_4_6 | (
    match_exuwbu_3_6 | (match_exuwbu_2_6 | (match_exuwbu_1_6 | match_exuwbu_0_6)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__out_7_ready = match_exuwbu_7_7 | (match_exuwbu_6_7 | (match_exuwbu_5_7 | (match_exuwbu_4_7 | (
    match_exuwbu_3_7 | (match_exuwbu_2_7 | (match_exuwbu_1_7 | match_exuwbu_0_7)))))); // @[Backend.scala 866:202 867:29]
  assign exu_io__flush = io_flush[1]; // @[Backend.scala 902:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[Backend.scala 933:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[Backend.scala 933:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Backend.scala 933:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[Backend.scala 932:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[Backend.scala 932:18]
  assign exu_io__memMMU_dmem_addr = io_memMMU_dmem_addr; // @[Backend.scala 932:18]
  assign exu__T_408 = _T_408_0;
  assign exu__T_137_0 = wbu__T_137_0;
  assign exu__T_140_0 = wbu__T_140_0;
  assign exu_io_in_0_valid = wbu_io_in_0_valid;
  assign exu_ismmio = ismmio;
  assign exu__WIRE_2_1 = wbu__WIRE_2_1;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu__T_136_0 = wbu__T_136_0;
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu__T_139_0 = wbu__T_139_0;
  assign exu_vmEnable = vmEnable;
  assign exu__T_407 = _T_407_0;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu__T_138_0 = wbu__T_138_0;
  assign exu__T_135_0 = wbu__T_135_0;
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io__in_0_valid = wbu_valid_0; // @[Backend.scala 842:24]
  assign wbu_io__in_0_bits_decode_cf_pc = wbu_bits_0_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_cf_redirect_target = wbu_bits_0_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_cf_redirect_valid = wbu_bits_0_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_cf_runahead_checkpoint_id = wbu_bits_0_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_ctrl_rfWen = wbu_bits_0_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_ctrl_rfDest = wbu_bits_0_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_pext_OV = wbu_bits_0_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_decode_InstNo = wbu_bits_0_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_0_bits_commits = wbu_bits_0_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_1_valid = wbu_valid_1; // @[Backend.scala 842:24]
  assign wbu_io__in_1_bits_decode_cf_pc = wbu_bits_1_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_cf_redirect_target = wbu_bits_1_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_cf_redirect_valid = wbu_bits_1_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_cf_runahead_checkpoint_id = wbu_bits_1_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_ctrl_rfWen = wbu_bits_1_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_ctrl_rfDest = wbu_bits_1_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_pext_OV = wbu_bits_1_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_decode_InstNo = wbu_bits_1_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_1_bits_commits = wbu_bits_1_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_2_valid = wbu_valid_2; // @[Backend.scala 842:24]
  assign wbu_io__in_2_bits_decode_cf_pc = wbu_bits_2_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_cf_redirect_target = wbu_bits_2_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_cf_redirect_valid = wbu_bits_2_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_cf_runahead_checkpoint_id = wbu_bits_2_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_ctrl_rfWen = wbu_bits_2_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_ctrl_rfDest = wbu_bits_2_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_pext_OV = wbu_bits_2_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_decode_InstNo = wbu_bits_2_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_2_bits_commits = wbu_bits_2_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_3_valid = wbu_valid_3; // @[Backend.scala 842:24]
  assign wbu_io__in_3_bits_decode_cf_pc = wbu_bits_3_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_cf_redirect_target = wbu_bits_3_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_cf_redirect_valid = wbu_bits_3_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_cf_runahead_checkpoint_id = wbu_bits_3_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_ctrl_rfWen = wbu_bits_3_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_ctrl_rfDest = wbu_bits_3_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_pext_OV = wbu_bits_3_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_decode_InstNo = wbu_bits_3_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_3_bits_commits = wbu_bits_3_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_4_valid = wbu_valid_4; // @[Backend.scala 842:24]
  assign wbu_io__in_4_bits_decode_cf_pc = wbu_bits_4_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_cf_redirect_target = wbu_bits_4_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_cf_redirect_valid = wbu_bits_4_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_cf_runahead_checkpoint_id = wbu_bits_4_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_ctrl_rfWen = wbu_bits_4_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_ctrl_rfDest = wbu_bits_4_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_pext_OV = wbu_bits_4_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_decode_InstNo = wbu_bits_4_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_4_bits_commits = wbu_bits_4_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_5_valid = wbu_valid_5; // @[Backend.scala 842:24]
  assign wbu_io__in_5_bits_decode_cf_pc = wbu_bits_5_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_cf_redirect_target = wbu_bits_5_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_cf_redirect_valid = wbu_bits_5_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_cf_runahead_checkpoint_id = wbu_bits_5_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_ctrl_rfWen = wbu_bits_5_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_ctrl_rfDest = wbu_bits_5_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_pext_OV = wbu_bits_5_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_decode_InstNo = wbu_bits_5_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_5_bits_commits = wbu_bits_5_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_6_valid = wbu_valid_6; // @[Backend.scala 842:24]
  assign wbu_io__in_6_bits_decode_cf_pc = wbu_bits_6_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_cf_redirect_target = wbu_bits_6_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_cf_redirect_valid = wbu_bits_6_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_cf_runahead_checkpoint_id = wbu_bits_6_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_ctrl_rfWen = wbu_bits_6_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_ctrl_rfDest = wbu_bits_6_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_pext_OV = wbu_bits_6_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_decode_InstNo = wbu_bits_6_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_6_bits_commits = wbu_bits_6_commits; // @[Backend.scala 841:23]
  assign wbu_io__in_7_valid = wbu_valid_7; // @[Backend.scala 842:24]
  assign wbu_io__in_7_bits_decode_cf_pc = wbu_bits_7_decode_cf_pc; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_cf_redirect_target = wbu_bits_7_decode_cf_redirect_target; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_cf_redirect_valid = wbu_bits_7_decode_cf_redirect_valid; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_cf_runahead_checkpoint_id = wbu_bits_7_decode_cf_runahead_checkpoint_id; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_ctrl_rfWen = wbu_bits_7_decode_ctrl_rfWen; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_ctrl_rfDest = wbu_bits_7_decode_ctrl_rfDest; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_pext_OV = wbu_bits_7_decode_pext_OV; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_decode_InstNo = wbu_bits_7_decode_InstNo; // @[Backend.scala 841:23]
  assign wbu_io__in_7_bits_commits = wbu_bits_7_commits; // @[Backend.scala 841:23]
  assign wbu_io__wb_rfSrc1_0 = isu_io_wb_rfSrc1_0; // @[Backend.scala 914:24]
  assign wbu_io__wb_rfSrc1_1 = isu_io_wb_rfSrc1_1; // @[Backend.scala 914:24]
  assign wbu_io__wb_rfSrc2_0 = isu_io_wb_rfSrc2_0; // @[Backend.scala 915:24]
  assign wbu_io__wb_rfSrc2_1 = isu_io_wb_rfSrc2_1; // @[Backend.scala 915:24]
  assign wbu_io__wb_rfSrc3_0 = isu_io_wb_rfSrc3_0; // @[Backend.scala 920:26]
  assign wbu_io__wb_rfSrc3_1 = isu_io_wb_rfSrc3_1; // @[Backend.scala 920:26]
  always @(posedge clock) begin
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_cf_instr <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_instr <= isu_io_out_1_bits_cf_instr; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_instr <= isu_io_out_0_bits_cf_instr; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_cf_pnpc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_pnpc <= isu_io_out_1_bits_cf_pnpc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_pnpc <= isu_io_out_0_bits_cf_pnpc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_cf_brIdx <= 4'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_brIdx <= isu_io_out_1_bits_cf_brIdx; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_brIdx <= isu_io_out_0_bits_cf_brIdx; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_data_imm <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_data_imm <= isu_io_out_1_bits_data_imm; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_data_imm <= isu_io_out_0_bits_data_imm; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_0_InstFlag <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_0) begin // @[Backend.scala 805:244]
      exu_bits_0_InstFlag <= isu_io_out_1_bits_InstFlag; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_0) begin // @[Backend.scala 805:244]
      exu_bits_0_InstFlag <= isu_io_out_0_bits_InstFlag; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_exceptionVec_1 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_exceptionVec_1 <= isu_io_out_1_bits_cf_exceptionVec_1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_exceptionVec_1 <= isu_io_out_0_bits_cf_exceptionVec_1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_exceptionVec_2 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_exceptionVec_2 <= isu_io_out_1_bits_cf_exceptionVec_2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_exceptionVec_2 <= isu_io_out_0_bits_cf_exceptionVec_2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_exceptionVec_12 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_exceptionVec_12 <= isu_io_out_1_bits_cf_exceptionVec_12; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_exceptionVec_12 <= isu_io_out_0_bits_cf_exceptionVec_12; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_0 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_0 <= isu_io_out_1_bits_cf_intrVec_0; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_0 <= isu_io_out_0_bits_cf_intrVec_0; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_1 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_1 <= isu_io_out_1_bits_cf_intrVec_1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_1 <= isu_io_out_0_bits_cf_intrVec_1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_2 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_2 <= isu_io_out_1_bits_cf_intrVec_2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_2 <= isu_io_out_0_bits_cf_intrVec_2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_3 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_3 <= isu_io_out_1_bits_cf_intrVec_3; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_3 <= isu_io_out_0_bits_cf_intrVec_3; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_4 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_4 <= isu_io_out_1_bits_cf_intrVec_4; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_4 <= isu_io_out_0_bits_cf_intrVec_4; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_5 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_5 <= isu_io_out_1_bits_cf_intrVec_5; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_5 <= isu_io_out_0_bits_cf_intrVec_5; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_6 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_6 <= isu_io_out_1_bits_cf_intrVec_6; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_6 <= isu_io_out_0_bits_cf_intrVec_6; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_7 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_7 <= isu_io_out_1_bits_cf_intrVec_7; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_7 <= isu_io_out_0_bits_cf_intrVec_7; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_8 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_8 <= isu_io_out_1_bits_cf_intrVec_8; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_8 <= isu_io_out_0_bits_cf_intrVec_8; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_9 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_9 <= isu_io_out_1_bits_cf_intrVec_9; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_9 <= isu_io_out_0_bits_cf_intrVec_9; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_10 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_10 <= isu_io_out_1_bits_cf_intrVec_10; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_10 <= isu_io_out_0_bits_cf_intrVec_10; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_intrVec_11 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_11 <= isu_io_out_1_bits_cf_intrVec_11; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_intrVec_11 <= isu_io_out_0_bits_cf_intrVec_11; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_crossPageIPFFix <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_crossPageIPFFix <= isu_io_out_1_bits_cf_crossPageIPFFix; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_crossPageIPFFix <= isu_io_out_0_bits_cf_crossPageIPFFix; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_ctrl_isMou <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_isMou <= isu_io_out_1_bits_ctrl_isMou; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_ctrl_isMou <= isu_io_out_0_bits_ctrl_isMou; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_1_InstFlag <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_1) begin // @[Backend.scala 805:244]
      exu_bits_1_InstFlag <= isu_io_out_1_bits_InstFlag; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_1) begin // @[Backend.scala 805:244]
      exu_bits_1_InstFlag <= isu_io_out_0_bits_InstFlag; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_cf_instr <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_instr <= isu_io_out_1_bits_cf_instr; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_instr <= isu_io_out_0_bits_cf_instr; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_cf_instrType <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_instrType <= isu_io_out_1_bits_cf_instrType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_cf_instrType <= isu_io_out_0_bits_cf_instrType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_ctrl_funct3 <= 3'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_funct3 <= isu_io_out_1_bits_ctrl_funct3; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_funct3 <= isu_io_out_0_bits_ctrl_funct3; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_ctrl_func24 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_func24 <= isu_io_out_1_bits_ctrl_func24; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_func24 <= isu_io_out_0_bits_ctrl_func24; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_ctrl_func23 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_func23 <= isu_io_out_1_bits_ctrl_func23; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_func23 <= isu_io_out_0_bits_ctrl_func23; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_data_src3 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_data_src3 <= isu_io_out_1_bits_data_src3; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_data_src3 <= isu_io_out_0_bits_data_src3; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_2_InstFlag <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_2) begin // @[Backend.scala 805:244]
      exu_bits_2_InstFlag <= isu_io_out_1_bits_InstFlag; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_2) begin // @[Backend.scala 805:244]
      exu_bits_2_InstFlag <= isu_io_out_0_bits_InstFlag; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_cf_instr <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_instr <= isu_io_out_1_bits_cf_instr; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_instr <= isu_io_out_0_bits_cf_instr; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_cf_instrType <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_instrType <= isu_io_out_1_bits_cf_instrType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_cf_instrType <= isu_io_out_0_bits_cf_instrType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_ctrl_funct3 <= 3'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_funct3 <= isu_io_out_1_bits_ctrl_funct3; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_funct3 <= isu_io_out_0_bits_ctrl_funct3; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_ctrl_func24 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_func24 <= isu_io_out_1_bits_ctrl_func24; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_func24 <= isu_io_out_0_bits_ctrl_func24; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_ctrl_func23 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_func23 <= isu_io_out_1_bits_ctrl_func23; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_func23 <= isu_io_out_0_bits_ctrl_func23; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_data_src3 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_data_src3 <= isu_io_out_1_bits_data_src3; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_data_src3 <= isu_io_out_0_bits_data_src3; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_3_InstFlag <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_3) begin // @[Backend.scala 805:244]
      exu_bits_3_InstFlag <= isu_io_out_1_bits_InstFlag; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_3) begin // @[Backend.scala 805:244]
      exu_bits_3_InstFlag <= isu_io_out_0_bits_InstFlag; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_instr <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_instr <= isu_io_out_1_bits_cf_instr; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_instr <= isu_io_out_0_bits_cf_instr; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_exceptionVec_1 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_exceptionVec_1 <= isu_io_out_1_bits_cf_exceptionVec_1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_exceptionVec_1 <= isu_io_out_0_bits_cf_exceptionVec_1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_exceptionVec_2 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_exceptionVec_2 <= isu_io_out_1_bits_cf_exceptionVec_2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_exceptionVec_2 <= isu_io_out_0_bits_cf_exceptionVec_2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_exceptionVec_12 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_exceptionVec_12 <= isu_io_out_1_bits_cf_exceptionVec_12; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_exceptionVec_12 <= isu_io_out_0_bits_cf_exceptionVec_12; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_0 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_0 <= isu_io_out_1_bits_cf_intrVec_0; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_0 <= isu_io_out_0_bits_cf_intrVec_0; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_1 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_1 <= isu_io_out_1_bits_cf_intrVec_1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_1 <= isu_io_out_0_bits_cf_intrVec_1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_2 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_2 <= isu_io_out_1_bits_cf_intrVec_2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_2 <= isu_io_out_0_bits_cf_intrVec_2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_3 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_3 <= isu_io_out_1_bits_cf_intrVec_3; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_3 <= isu_io_out_0_bits_cf_intrVec_3; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_4 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_4 <= isu_io_out_1_bits_cf_intrVec_4; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_4 <= isu_io_out_0_bits_cf_intrVec_4; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_5 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_5 <= isu_io_out_1_bits_cf_intrVec_5; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_5 <= isu_io_out_0_bits_cf_intrVec_5; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_6 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_6 <= isu_io_out_1_bits_cf_intrVec_6; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_6 <= isu_io_out_0_bits_cf_intrVec_6; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_7 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_7 <= isu_io_out_1_bits_cf_intrVec_7; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_7 <= isu_io_out_0_bits_cf_intrVec_7; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_8 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_8 <= isu_io_out_1_bits_cf_intrVec_8; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_8 <= isu_io_out_0_bits_cf_intrVec_8; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_9 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_9 <= isu_io_out_1_bits_cf_intrVec_9; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_9 <= isu_io_out_0_bits_cf_intrVec_9; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_10 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_10 <= isu_io_out_1_bits_cf_intrVec_10; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_10 <= isu_io_out_0_bits_cf_intrVec_10; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_intrVec_11 <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_11 <= isu_io_out_1_bits_cf_intrVec_11; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_intrVec_11 <= isu_io_out_0_bits_cf_intrVec_11; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_crossPageIPFFix <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_crossPageIPFFix <= isu_io_out_1_bits_cf_crossPageIPFFix; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_crossPageIPFFix <= isu_io_out_0_bits_cf_crossPageIPFFix; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_ctrl_isMou <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_isMou <= isu_io_out_1_bits_ctrl_isMou; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_ctrl_isMou <= isu_io_out_0_bits_ctrl_isMou; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_data_imm <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_data_imm <= isu_io_out_1_bits_data_imm; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_data_imm <= isu_io_out_0_bits_data_imm; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_4_InstFlag <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_4) begin // @[Backend.scala 805:244]
      exu_bits_4_InstFlag <= isu_io_out_1_bits_InstFlag; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_4) begin // @[Backend.scala 805:244]
      exu_bits_4_InstFlag <= isu_io_out_0_bits_InstFlag; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_5_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_5) begin // @[Backend.scala 805:244]
      exu_bits_5_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_5) begin // @[Backend.scala 805:244]
      exu_bits_5_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_cf_instr <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_instr <= isu_io_out_1_bits_cf_instr; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_instr <= isu_io_out_0_bits_cf_instr; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_cf_pnpc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_pnpc <= isu_io_out_1_bits_cf_pnpc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_pnpc <= isu_io_out_0_bits_cf_pnpc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_cf_brIdx <= 4'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_brIdx <= isu_io_out_1_bits_cf_brIdx; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_brIdx <= isu_io_out_0_bits_cf_brIdx; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_data_imm <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_data_imm <= isu_io_out_1_bits_data_imm; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_data_imm <= isu_io_out_0_bits_data_imm; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_6_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_6) begin // @[Backend.scala 805:244]
      exu_bits_6_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_6) begin // @[Backend.scala 805:244]
      exu_bits_6_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_cf_instr <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_instr <= isu_io_out_1_bits_cf_instr; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_instr <= isu_io_out_0_bits_cf_instr; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_cf_pc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_pc <= isu_io_out_1_bits_cf_pc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_pc <= isu_io_out_0_bits_cf_pc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_cf_pnpc <= 39'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_pnpc <= isu_io_out_1_bits_cf_pnpc; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_pnpc <= isu_io_out_0_bits_cf_pnpc; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_cf_brIdx <= 4'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_brIdx <= isu_io_out_1_bits_cf_brIdx; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_brIdx <= isu_io_out_0_bits_cf_brIdx; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_runahead_checkpoint_id <= isu_io_out_1_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_cf_runahead_checkpoint_id <= isu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_ctrl_fuOpType <= 7'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_ctrl_fuOpType <= isu_io_out_1_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_ctrl_fuOpType <= isu_io_out_0_bits_ctrl_fuOpType; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_ctrl_rfWen <= 1'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_ctrl_rfWen <= isu_io_out_1_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_ctrl_rfWen <= isu_io_out_0_bits_ctrl_rfWen; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_ctrl_rfDest <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_ctrl_rfDest <= isu_io_out_1_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_ctrl_rfDest <= isu_io_out_0_bits_ctrl_rfDest; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_data_src1 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_data_src1 <= isu_io_out_1_bits_data_src1; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_data_src1 <= isu_io_out_0_bits_data_src1; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_data_src2 <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_data_src2 <= isu_io_out_1_bits_data_src2; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_data_src2 <= isu_io_out_0_bits_data_src2; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_data_imm <= 64'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_data_imm <= isu_io_out_1_bits_data_imm; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_data_imm <= isu_io_out_0_bits_data_imm; // @[Backend.scala 808:28]
    end
    if (reset) begin // @[Backend.scala 732:30]
      exu_bits_7_InstNo <= 5'h0; // @[Backend.scala 732:30]
    end else if (match_operaotr_1_7) begin // @[Backend.scala 805:244]
      exu_bits_7_InstNo <= isu_io_out_1_bits_InstNo; // @[Backend.scala 808:28]
    end else if (match_operaotr_0_7) begin // @[Backend.scala 805:244]
      exu_bits_7_InstNo <= isu_io_out_0_bits_InstNo; // @[Backend.scala 808:28]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_0 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_0 <= exu_valid_next_0; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_1 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_1 <= exu_valid_next_1; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_2 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_2 <= exu_valid_next_2; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_3 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_3 <= exu_valid_next_3; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_4 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_4 <= exu_valid_next_4; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_5 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_5 <= exu_valid_next_5; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_6 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_6 <= exu_valid_next_6; // @[Backend.scala 823:15]
    end
    if (reset | io_flush[0]) begin // @[Backend.scala 820:36]
      exu_valid_7 <= 1'h0; // @[Backend.scala 821:47]
    end else begin
      exu_valid_7 <= exu_valid_next_7; // @[Backend.scala 823:15]
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_cf_pc <= _GEN_1484;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_cf_redirect_target <= _GEN_1482;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_cf_redirect_valid <= _GEN_1480;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_cf_runahead_checkpoint_id <= _GEN_1448;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_ctrl_rfWen <= _GEN_1435;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_ctrl_rfDest <= _GEN_1434;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_pext_OV <= _GEN_1422;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_decode_InstNo <= _GEN_1421;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_0_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_0_7) begin // @[Backend.scala 866:202]
      wbu_bits_0_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_6) begin // @[Backend.scala 866:202]
      wbu_bits_0_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_0_5) begin // @[Backend.scala 866:202]
      wbu_bits_0_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_0_commits <= _GEN_1417;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_cf_pc <= _GEN_2060;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_cf_redirect_target <= _GEN_2058;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_cf_redirect_valid <= _GEN_2056;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_cf_runahead_checkpoint_id <= _GEN_2024;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_ctrl_rfWen <= _GEN_2011;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_ctrl_rfDest <= _GEN_2010;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_pext_OV <= _GEN_1998;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_decode_InstNo <= _GEN_1997;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_1_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_1_7) begin // @[Backend.scala 866:202]
      wbu_bits_1_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_6) begin // @[Backend.scala 866:202]
      wbu_bits_1_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_1_5) begin // @[Backend.scala 866:202]
      wbu_bits_1_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_1_commits <= _GEN_1993;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_cf_pc <= _GEN_2636;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_cf_redirect_target <= _GEN_2634;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_cf_redirect_valid <= _GEN_2632;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_cf_runahead_checkpoint_id <= _GEN_2600;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_ctrl_rfWen <= _GEN_2587;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_ctrl_rfDest <= _GEN_2586;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_pext_OV <= _GEN_2574;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_decode_InstNo <= _GEN_2573;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_2_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_2_7) begin // @[Backend.scala 866:202]
      wbu_bits_2_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_6) begin // @[Backend.scala 866:202]
      wbu_bits_2_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_2_5) begin // @[Backend.scala 866:202]
      wbu_bits_2_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_2_commits <= _GEN_2569;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_cf_pc <= _GEN_3212;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_cf_redirect_target <= _GEN_3210;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_cf_redirect_valid <= _GEN_3208;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_cf_runahead_checkpoint_id <= _GEN_3176;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_ctrl_rfWen <= _GEN_3163;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_ctrl_rfDest <= _GEN_3162;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_pext_OV <= _GEN_3150;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_decode_InstNo <= _GEN_3149;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_3_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_3_7) begin // @[Backend.scala 866:202]
      wbu_bits_3_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_6) begin // @[Backend.scala 866:202]
      wbu_bits_3_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_3_5) begin // @[Backend.scala 866:202]
      wbu_bits_3_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_3_commits <= _GEN_3145;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_cf_pc <= _GEN_3788;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_cf_redirect_target <= _GEN_3786;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_cf_redirect_valid <= _GEN_3784;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_cf_runahead_checkpoint_id <= _GEN_3752;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_ctrl_rfWen <= _GEN_3739;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_ctrl_rfDest <= _GEN_3738;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_pext_OV <= _GEN_3726;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_decode_InstNo <= _GEN_3725;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_4_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_4_7) begin // @[Backend.scala 866:202]
      wbu_bits_4_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_6) begin // @[Backend.scala 866:202]
      wbu_bits_4_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_4_5) begin // @[Backend.scala 866:202]
      wbu_bits_4_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_4_commits <= _GEN_3721;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_cf_pc <= _GEN_4364;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_cf_redirect_target <= _GEN_4362;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_cf_redirect_valid <= _GEN_4360;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_cf_runahead_checkpoint_id <= _GEN_4328;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_ctrl_rfWen <= _GEN_4315;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_ctrl_rfDest <= _GEN_4314;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_pext_OV <= _GEN_4302;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_decode_InstNo <= _GEN_4301;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_5_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_5_7) begin // @[Backend.scala 866:202]
      wbu_bits_5_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_6) begin // @[Backend.scala 866:202]
      wbu_bits_5_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_5_5) begin // @[Backend.scala 866:202]
      wbu_bits_5_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_5_commits <= _GEN_4297;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_cf_pc <= _GEN_4940;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_cf_redirect_target <= _GEN_4938;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_cf_redirect_valid <= _GEN_4936;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_cf_runahead_checkpoint_id <= _GEN_4904;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_ctrl_rfWen <= _GEN_4891;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_ctrl_rfDest <= _GEN_4890;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_pext_OV <= _GEN_4878;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_decode_InstNo <= _GEN_4877;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_6_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_6_7) begin // @[Backend.scala 866:202]
      wbu_bits_6_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_6) begin // @[Backend.scala 866:202]
      wbu_bits_6_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_6_5) begin // @[Backend.scala 866:202]
      wbu_bits_6_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_6_commits <= _GEN_4873;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_cf_pc <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_pc <= exu_io__out_7_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_pc <= exu_io__out_6_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_pc <= exu_io__out_5_bits_decode_cf_pc; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_cf_pc <= _GEN_5516;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_redirect_target <= exu_io__out_7_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_redirect_target <= exu_io__out_6_bits_decode_cf_redirect_target; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_redirect_target <= 39'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_cf_redirect_target <= _GEN_5514;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_redirect_valid <= exu_io__out_7_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_redirect_valid <= exu_io__out_6_bits_decode_cf_redirect_valid; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_redirect_valid <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_cf_redirect_valid <= _GEN_5512;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_cf_runahead_checkpoint_id <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_runahead_checkpoint_id <= exu_io__out_7_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_runahead_checkpoint_id <= exu_io__out_6_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_cf_runahead_checkpoint_id <= exu_io__out_5_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_cf_runahead_checkpoint_id <= _GEN_5480;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_ctrl_rfWen <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_ctrl_rfWen <= exu_io__out_7_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_ctrl_rfWen <= exu_io__out_6_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_ctrl_rfWen <= exu_io__out_5_bits_decode_ctrl_rfWen; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_ctrl_rfWen <= _GEN_5467;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_ctrl_rfDest <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_ctrl_rfDest <= exu_io__out_7_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_ctrl_rfDest <= exu_io__out_6_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_ctrl_rfDest <= exu_io__out_5_bits_decode_ctrl_rfDest; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_ctrl_rfDest <= _GEN_5466;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_pext_OV <= 1'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_pext_OV <= 1'h0; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_pext_OV <= _GEN_5454;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_decode_InstNo <= 5'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_InstNo <= exu_io__out_7_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_InstNo <= exu_io__out_6_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_decode_InstNo <= exu_io__out_5_bits_decode_InstNo; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_decode_InstNo <= _GEN_5453;
    end
    if (reset) begin // @[Backend.scala 833:30]
      wbu_bits_7_commits <= 64'h0; // @[Backend.scala 833:30]
    end else if (match_exuwbu_7_7) begin // @[Backend.scala 866:202]
      wbu_bits_7_commits <= exu_io__out_7_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_6) begin // @[Backend.scala 866:202]
      wbu_bits_7_commits <= exu_io__out_6_bits_commits; // @[Backend.scala 868:26]
    end else if (match_exuwbu_7_5) begin // @[Backend.scala 866:202]
      wbu_bits_7_commits <= exu_io__out_5_bits_commits; // @[Backend.scala 868:26]
    end else begin
      wbu_bits_7_commits <= _GEN_5449;
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_0 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_0 <= wbu_valid_next_0; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_1 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_1 <= wbu_valid_next_1; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_2 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_2 <= wbu_valid_next_2; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_3 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_3 <= wbu_valid_next_3; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_4 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_4 <= wbu_valid_next_4; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_5 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_5 <= wbu_valid_next_5; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_6 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_6 <= wbu_valid_next_6; // @[Backend.scala 888:14]
    end
    if (reset) begin // @[Backend.scala 885:21]
      wbu_valid_7 <= 1'h0; // @[Backend.scala 886:47]
    end else begin
      wbu_valid_7 <= wbu_valid_next_7; // @[Backend.scala 888:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  exu_bits_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  exu_bits_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  exu_bits_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  exu_bits_0_cf_brIdx = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  exu_bits_0_cf_runahead_checkpoint_id = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  exu_bits_0_ctrl_fuOpType = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  exu_bits_0_ctrl_rfWen = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exu_bits_0_ctrl_rfDest = _RAND_7[4:0];
  _RAND_8 = {2{`RANDOM}};
  exu_bits_0_data_src1 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  exu_bits_0_data_src2 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  exu_bits_0_data_imm = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  exu_bits_0_InstNo = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  exu_bits_0_InstFlag = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  exu_bits_1_cf_pc = _RAND_13[38:0];
  _RAND_14 = {1{`RANDOM}};
  exu_bits_1_cf_exceptionVec_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exu_bits_1_cf_exceptionVec_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  exu_bits_1_cf_exceptionVec_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_3 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_4 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_5 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_6 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_7 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_8 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_9 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_10 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  exu_bits_1_cf_intrVec_11 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  exu_bits_1_cf_crossPageIPFFix = _RAND_29[0:0];
  _RAND_30 = {2{`RANDOM}};
  exu_bits_1_cf_runahead_checkpoint_id = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  exu_bits_1_ctrl_fuOpType = _RAND_31[6:0];
  _RAND_32 = {1{`RANDOM}};
  exu_bits_1_ctrl_rfWen = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  exu_bits_1_ctrl_rfDest = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  exu_bits_1_ctrl_isMou = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  exu_bits_1_data_src1 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  exu_bits_1_data_src2 = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  exu_bits_1_InstNo = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  exu_bits_1_InstFlag = _RAND_38[0:0];
  _RAND_39 = {2{`RANDOM}};
  exu_bits_2_cf_instr = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  exu_bits_2_cf_pc = _RAND_40[38:0];
  _RAND_41 = {2{`RANDOM}};
  exu_bits_2_cf_runahead_checkpoint_id = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  exu_bits_2_cf_instrType = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  exu_bits_2_ctrl_fuOpType = _RAND_43[6:0];
  _RAND_44 = {1{`RANDOM}};
  exu_bits_2_ctrl_funct3 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  exu_bits_2_ctrl_func24 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  exu_bits_2_ctrl_func23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  exu_bits_2_ctrl_rfWen = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  exu_bits_2_ctrl_rfDest = _RAND_48[4:0];
  _RAND_49 = {2{`RANDOM}};
  exu_bits_2_data_src1 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  exu_bits_2_data_src2 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  exu_bits_2_data_src3 = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  exu_bits_2_InstNo = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  exu_bits_2_InstFlag = _RAND_53[0:0];
  _RAND_54 = {2{`RANDOM}};
  exu_bits_3_cf_instr = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  exu_bits_3_cf_pc = _RAND_55[38:0];
  _RAND_56 = {2{`RANDOM}};
  exu_bits_3_cf_runahead_checkpoint_id = _RAND_56[63:0];
  _RAND_57 = {1{`RANDOM}};
  exu_bits_3_cf_instrType = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  exu_bits_3_ctrl_fuOpType = _RAND_58[6:0];
  _RAND_59 = {1{`RANDOM}};
  exu_bits_3_ctrl_funct3 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  exu_bits_3_ctrl_func24 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  exu_bits_3_ctrl_func23 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  exu_bits_3_ctrl_rfWen = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  exu_bits_3_ctrl_rfDest = _RAND_63[4:0];
  _RAND_64 = {2{`RANDOM}};
  exu_bits_3_data_src1 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  exu_bits_3_data_src2 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  exu_bits_3_data_src3 = _RAND_66[63:0];
  _RAND_67 = {1{`RANDOM}};
  exu_bits_3_InstNo = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  exu_bits_3_InstFlag = _RAND_68[0:0];
  _RAND_69 = {2{`RANDOM}};
  exu_bits_4_cf_instr = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  exu_bits_4_cf_pc = _RAND_70[38:0];
  _RAND_71 = {1{`RANDOM}};
  exu_bits_4_cf_exceptionVec_1 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  exu_bits_4_cf_exceptionVec_2 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  exu_bits_4_cf_exceptionVec_12 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_3 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_4 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_5 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_6 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_8 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_9 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_10 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  exu_bits_4_cf_intrVec_11 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  exu_bits_4_cf_crossPageIPFFix = _RAND_86[0:0];
  _RAND_87 = {2{`RANDOM}};
  exu_bits_4_cf_runahead_checkpoint_id = _RAND_87[63:0];
  _RAND_88 = {1{`RANDOM}};
  exu_bits_4_ctrl_fuOpType = _RAND_88[6:0];
  _RAND_89 = {1{`RANDOM}};
  exu_bits_4_ctrl_rfWen = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  exu_bits_4_ctrl_rfDest = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  exu_bits_4_ctrl_isMou = _RAND_91[0:0];
  _RAND_92 = {2{`RANDOM}};
  exu_bits_4_data_src1 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  exu_bits_4_data_src2 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  exu_bits_4_data_imm = _RAND_94[63:0];
  _RAND_95 = {1{`RANDOM}};
  exu_bits_4_InstNo = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  exu_bits_4_InstFlag = _RAND_96[0:0];
  _RAND_97 = {2{`RANDOM}};
  exu_bits_5_cf_pc = _RAND_97[38:0];
  _RAND_98 = {2{`RANDOM}};
  exu_bits_5_cf_runahead_checkpoint_id = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  exu_bits_5_ctrl_fuOpType = _RAND_99[6:0];
  _RAND_100 = {1{`RANDOM}};
  exu_bits_5_ctrl_rfWen = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  exu_bits_5_ctrl_rfDest = _RAND_101[4:0];
  _RAND_102 = {2{`RANDOM}};
  exu_bits_5_data_src1 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  exu_bits_5_data_src2 = _RAND_103[63:0];
  _RAND_104 = {1{`RANDOM}};
  exu_bits_5_InstNo = _RAND_104[4:0];
  _RAND_105 = {2{`RANDOM}};
  exu_bits_6_cf_instr = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  exu_bits_6_cf_pc = _RAND_106[38:0];
  _RAND_107 = {2{`RANDOM}};
  exu_bits_6_cf_pnpc = _RAND_107[38:0];
  _RAND_108 = {1{`RANDOM}};
  exu_bits_6_cf_brIdx = _RAND_108[3:0];
  _RAND_109 = {2{`RANDOM}};
  exu_bits_6_cf_runahead_checkpoint_id = _RAND_109[63:0];
  _RAND_110 = {1{`RANDOM}};
  exu_bits_6_ctrl_fuOpType = _RAND_110[6:0];
  _RAND_111 = {1{`RANDOM}};
  exu_bits_6_ctrl_rfWen = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  exu_bits_6_ctrl_rfDest = _RAND_112[4:0];
  _RAND_113 = {2{`RANDOM}};
  exu_bits_6_data_src1 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  exu_bits_6_data_src2 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  exu_bits_6_data_imm = _RAND_115[63:0];
  _RAND_116 = {1{`RANDOM}};
  exu_bits_6_InstNo = _RAND_116[4:0];
  _RAND_117 = {2{`RANDOM}};
  exu_bits_7_cf_instr = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  exu_bits_7_cf_pc = _RAND_118[38:0];
  _RAND_119 = {2{`RANDOM}};
  exu_bits_7_cf_pnpc = _RAND_119[38:0];
  _RAND_120 = {1{`RANDOM}};
  exu_bits_7_cf_brIdx = _RAND_120[3:0];
  _RAND_121 = {2{`RANDOM}};
  exu_bits_7_cf_runahead_checkpoint_id = _RAND_121[63:0];
  _RAND_122 = {1{`RANDOM}};
  exu_bits_7_ctrl_fuOpType = _RAND_122[6:0];
  _RAND_123 = {1{`RANDOM}};
  exu_bits_7_ctrl_rfWen = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  exu_bits_7_ctrl_rfDest = _RAND_124[4:0];
  _RAND_125 = {2{`RANDOM}};
  exu_bits_7_data_src1 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  exu_bits_7_data_src2 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  exu_bits_7_data_imm = _RAND_127[63:0];
  _RAND_128 = {1{`RANDOM}};
  exu_bits_7_InstNo = _RAND_128[4:0];
  _RAND_129 = {1{`RANDOM}};
  exu_valid_0 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  exu_valid_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  exu_valid_2 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  exu_valid_3 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  exu_valid_4 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  exu_valid_5 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  exu_valid_6 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  exu_valid_7 = _RAND_136[0:0];
  _RAND_137 = {2{`RANDOM}};
  wbu_bits_0_decode_cf_pc = _RAND_137[38:0];
  _RAND_138 = {2{`RANDOM}};
  wbu_bits_0_decode_cf_redirect_target = _RAND_138[38:0];
  _RAND_139 = {1{`RANDOM}};
  wbu_bits_0_decode_cf_redirect_valid = _RAND_139[0:0];
  _RAND_140 = {2{`RANDOM}};
  wbu_bits_0_decode_cf_runahead_checkpoint_id = _RAND_140[63:0];
  _RAND_141 = {1{`RANDOM}};
  wbu_bits_0_decode_ctrl_rfWen = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  wbu_bits_0_decode_ctrl_rfDest = _RAND_142[4:0];
  _RAND_143 = {1{`RANDOM}};
  wbu_bits_0_decode_pext_OV = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  wbu_bits_0_decode_InstNo = _RAND_144[4:0];
  _RAND_145 = {2{`RANDOM}};
  wbu_bits_0_commits = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  wbu_bits_1_decode_cf_pc = _RAND_146[38:0];
  _RAND_147 = {2{`RANDOM}};
  wbu_bits_1_decode_cf_redirect_target = _RAND_147[38:0];
  _RAND_148 = {1{`RANDOM}};
  wbu_bits_1_decode_cf_redirect_valid = _RAND_148[0:0];
  _RAND_149 = {2{`RANDOM}};
  wbu_bits_1_decode_cf_runahead_checkpoint_id = _RAND_149[63:0];
  _RAND_150 = {1{`RANDOM}};
  wbu_bits_1_decode_ctrl_rfWen = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  wbu_bits_1_decode_ctrl_rfDest = _RAND_151[4:0];
  _RAND_152 = {1{`RANDOM}};
  wbu_bits_1_decode_pext_OV = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  wbu_bits_1_decode_InstNo = _RAND_153[4:0];
  _RAND_154 = {2{`RANDOM}};
  wbu_bits_1_commits = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  wbu_bits_2_decode_cf_pc = _RAND_155[38:0];
  _RAND_156 = {2{`RANDOM}};
  wbu_bits_2_decode_cf_redirect_target = _RAND_156[38:0];
  _RAND_157 = {1{`RANDOM}};
  wbu_bits_2_decode_cf_redirect_valid = _RAND_157[0:0];
  _RAND_158 = {2{`RANDOM}};
  wbu_bits_2_decode_cf_runahead_checkpoint_id = _RAND_158[63:0];
  _RAND_159 = {1{`RANDOM}};
  wbu_bits_2_decode_ctrl_rfWen = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  wbu_bits_2_decode_ctrl_rfDest = _RAND_160[4:0];
  _RAND_161 = {1{`RANDOM}};
  wbu_bits_2_decode_pext_OV = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  wbu_bits_2_decode_InstNo = _RAND_162[4:0];
  _RAND_163 = {2{`RANDOM}};
  wbu_bits_2_commits = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  wbu_bits_3_decode_cf_pc = _RAND_164[38:0];
  _RAND_165 = {2{`RANDOM}};
  wbu_bits_3_decode_cf_redirect_target = _RAND_165[38:0];
  _RAND_166 = {1{`RANDOM}};
  wbu_bits_3_decode_cf_redirect_valid = _RAND_166[0:0];
  _RAND_167 = {2{`RANDOM}};
  wbu_bits_3_decode_cf_runahead_checkpoint_id = _RAND_167[63:0];
  _RAND_168 = {1{`RANDOM}};
  wbu_bits_3_decode_ctrl_rfWen = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  wbu_bits_3_decode_ctrl_rfDest = _RAND_169[4:0];
  _RAND_170 = {1{`RANDOM}};
  wbu_bits_3_decode_pext_OV = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  wbu_bits_3_decode_InstNo = _RAND_171[4:0];
  _RAND_172 = {2{`RANDOM}};
  wbu_bits_3_commits = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  wbu_bits_4_decode_cf_pc = _RAND_173[38:0];
  _RAND_174 = {2{`RANDOM}};
  wbu_bits_4_decode_cf_redirect_target = _RAND_174[38:0];
  _RAND_175 = {1{`RANDOM}};
  wbu_bits_4_decode_cf_redirect_valid = _RAND_175[0:0];
  _RAND_176 = {2{`RANDOM}};
  wbu_bits_4_decode_cf_runahead_checkpoint_id = _RAND_176[63:0];
  _RAND_177 = {1{`RANDOM}};
  wbu_bits_4_decode_ctrl_rfWen = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  wbu_bits_4_decode_ctrl_rfDest = _RAND_178[4:0];
  _RAND_179 = {1{`RANDOM}};
  wbu_bits_4_decode_pext_OV = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  wbu_bits_4_decode_InstNo = _RAND_180[4:0];
  _RAND_181 = {2{`RANDOM}};
  wbu_bits_4_commits = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  wbu_bits_5_decode_cf_pc = _RAND_182[38:0];
  _RAND_183 = {2{`RANDOM}};
  wbu_bits_5_decode_cf_redirect_target = _RAND_183[38:0];
  _RAND_184 = {1{`RANDOM}};
  wbu_bits_5_decode_cf_redirect_valid = _RAND_184[0:0];
  _RAND_185 = {2{`RANDOM}};
  wbu_bits_5_decode_cf_runahead_checkpoint_id = _RAND_185[63:0];
  _RAND_186 = {1{`RANDOM}};
  wbu_bits_5_decode_ctrl_rfWen = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  wbu_bits_5_decode_ctrl_rfDest = _RAND_187[4:0];
  _RAND_188 = {1{`RANDOM}};
  wbu_bits_5_decode_pext_OV = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  wbu_bits_5_decode_InstNo = _RAND_189[4:0];
  _RAND_190 = {2{`RANDOM}};
  wbu_bits_5_commits = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  wbu_bits_6_decode_cf_pc = _RAND_191[38:0];
  _RAND_192 = {2{`RANDOM}};
  wbu_bits_6_decode_cf_redirect_target = _RAND_192[38:0];
  _RAND_193 = {1{`RANDOM}};
  wbu_bits_6_decode_cf_redirect_valid = _RAND_193[0:0];
  _RAND_194 = {2{`RANDOM}};
  wbu_bits_6_decode_cf_runahead_checkpoint_id = _RAND_194[63:0];
  _RAND_195 = {1{`RANDOM}};
  wbu_bits_6_decode_ctrl_rfWen = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  wbu_bits_6_decode_ctrl_rfDest = _RAND_196[4:0];
  _RAND_197 = {1{`RANDOM}};
  wbu_bits_6_decode_pext_OV = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  wbu_bits_6_decode_InstNo = _RAND_198[4:0];
  _RAND_199 = {2{`RANDOM}};
  wbu_bits_6_commits = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  wbu_bits_7_decode_cf_pc = _RAND_200[38:0];
  _RAND_201 = {2{`RANDOM}};
  wbu_bits_7_decode_cf_redirect_target = _RAND_201[38:0];
  _RAND_202 = {1{`RANDOM}};
  wbu_bits_7_decode_cf_redirect_valid = _RAND_202[0:0];
  _RAND_203 = {2{`RANDOM}};
  wbu_bits_7_decode_cf_runahead_checkpoint_id = _RAND_203[63:0];
  _RAND_204 = {1{`RANDOM}};
  wbu_bits_7_decode_ctrl_rfWen = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  wbu_bits_7_decode_ctrl_rfDest = _RAND_205[4:0];
  _RAND_206 = {1{`RANDOM}};
  wbu_bits_7_decode_pext_OV = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  wbu_bits_7_decode_InstNo = _RAND_207[4:0];
  _RAND_208 = {2{`RANDOM}};
  wbu_bits_7_commits = _RAND_208[63:0];
  _RAND_209 = {1{`RANDOM}};
  wbu_valid_0 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  wbu_valid_1 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  wbu_valid_2 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  wbu_valid_3 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  wbu_valid_4 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  wbu_valid_5 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  wbu_valid_6 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  wbu_valid_7 = _RAND_216[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] value; // @[Counter.scala 60:40]
  reg  lockIdx; // @[Arbiter.scala 46:22]
  wire  locked = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire  choice = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 88:{27,36}]
  wire  _T_2 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[Arbiter.scala 57:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : io_in_0_bits_size; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : io_in_0_bits_wmask; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:{15,15}]
  assign io_chosen = locked ? lockIdx : choice; // @[Arbiter.scala 40:13 55:{19,31}]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      lockIdx <= io_chosen; // @[Arbiter.scala 51:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [2:0]  io_in_1_req_bits_size,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [7:0]  io_in_1_req_bits_wmask,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 95:24]
  wire  inputArb_reset; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[Crossbar.scala 95:24]
  reg [1:0] state; // @[Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  reg  inflightSrc; // @[Crossbar.scala 99:28]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 103:47]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_25 | _T_26 ? 2'h2 : state; // @[Crossbar.scala 118:{80,88} 92:22]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [1:0] _GEN_9 = _T_29 ? 2'h0 : state; // @[Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter inputArb ( // @[Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 106:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 92:22]
      state <= 2'h0; // @[Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[Crossbar.scala 113:18]
      if (_T_19) begin // @[Crossbar.scala 115:29]
        if (_T_4) begin // @[Crossbar.scala 117:38]
          state <= 2'h1; // @[Crossbar.scala 117:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[Crossbar.scala 113:18]
      if (_T_29 & _T_30) begin // @[Crossbar.scala 121:82]
        state <= 2'h0; // @[Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[Crossbar.scala 113:18]
      state <= _GEN_9;
    end
    if (reset) begin // @[Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[Crossbar.scala 113:18]
      if (_T_19) begin // @[Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Crossbar.scala 98:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [3:0]  io_in_1_bits_cmd,
  input  [63:0] io_in_1_bits_wdata,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [3:0]  io_in_2_bits_cmd,
  input  [63:0] io_in_2_bits_wdata,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [2:0]  io_in_3_bits_size,
  input  [3:0]  io_in_3_bits_cmd,
  input  [7:0]  io_in_3_bits_wmask,
  input  [63:0] io_in_3_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 41:{16,16}]
  wire [63:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:{15,15}]
  wire [63:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_5; // @[Arbiter.scala 42:{15,15}]
  wire [7:0] _GEN_9 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[Arbiter.scala 42:{15,15}]
  wire [7:0] _GEN_10 = 2'h2 == io_chosen ? 8'hff : _GEN_9; // @[Arbiter.scala 42:{15,15}]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:{15,15}]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_13; // @[Arbiter.scala 42:{15,15}]
  wire [2:0] _GEN_17 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[Arbiter.scala 42:{15,15}]
  wire [2:0] _GEN_18 = 2'h2 == io_chosen ? 3'h3 : _GEN_17; // @[Arbiter.scala 42:{15,15}]
  wire [31:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:{15,15}]
  wire [31:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_21; // @[Arbiter.scala 42:{15,15}]
  reg [2:0] value; // @[Counter.scala 60:40]
  reg [1:0] lockIdx; // @[Arbiter.scala 46:22]
  wire  locked = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [1:0] _GEN_27 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 88:{27,36}]
  wire [1:0] _GEN_28 = io_in_1_valid ? 2'h1 : _GEN_27; // @[Arbiter.scala 88:{27,36}]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _GEN_28; // @[Arbiter.scala 88:{27,36}]
  wire  _T_4 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_5 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 31:78]
  wire  _T_6 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 31:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx == 2'h1 : _T_4; // @[Arbiter.scala 57:22]
  wire  _io_in_2_ready_T_1 = locked ? lockIdx == 2'h2 : _T_5; // @[Arbiter.scala 57:22]
  wire  _io_in_3_ready_T_1 = locked ? lockIdx == 2'h3 : _T_6; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_2_ready = _io_in_2_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_3_ready = _io_in_3_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 41:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_22; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_18; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_14; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_10; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_6; // @[Arbiter.scala 42:{15,15}]
  assign io_chosen = locked ? lockIdx : choice; // @[Arbiter.scala 40:13 55:{19,31}]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      lockIdx <= io_chosen; // @[Arbiter.scala 51:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input  [3:0]  io_in_2_req_bits_cmd,
  input  [63:0] io_in_2_req_bits_wdata,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input  [2:0]  io_in_3_req_bits_size,
  input  [3:0]  io_in_3_req_bits_cmd,
  input  [7:0]  io_in_3_req_bits_wmask,
  input  [63:0] io_in_3_req_bits_wdata,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [3:0]  io_in_3_resp_bits_cmd,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 95:24]
  wire  inputArb_reset; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_2_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_2_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_3_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_in_3_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 95:24]
  wire [1:0] inputArb_io_chosen; // @[Crossbar.scala 95:24]
  reg [1:0] state; // @[Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  reg [1:0] inflightSrc; // @[Crossbar.scala 99:28]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 103:47]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_25 | _T_26 ? 2'h2 : state; // @[Crossbar.scala 118:{80,88} 92:22]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [1:0] _GEN_13 = _T_29 ? 2'h0 : state; // @[Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter_1 inputArb ( // @[Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 96:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 96:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 106:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[Crossbar.scala 96:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 109:{13,13} 107:26]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 106:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[Crossbar.scala 96:68]
  assign io_in_3_resp_valid = 2'h3 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 109:{13,13} 107:26]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 106:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : 1'h1; // @[Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 92:22]
      state <= 2'h0; // @[Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[Crossbar.scala 113:18]
      if (_T_19) begin // @[Crossbar.scala 115:29]
        if (_T_4) begin // @[Crossbar.scala 117:38]
          state <= 2'h1; // @[Crossbar.scala 117:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (2'h1 == state) begin // @[Crossbar.scala 113:18]
      if (_T_29 & _T_30) begin // @[Crossbar.scala 121:82]
        state <= 2'h0; // @[Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[Crossbar.scala 113:18]
      state <= _GEN_13;
    end
    if (reset) begin // @[Crossbar.scala 99:28]
      inflightSrc <= 2'h0; // @[Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[Crossbar.scala 113:18]
      if (_T_19) begin // @[Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Crossbar.scala 98:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SIMD_TLBEXEC(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_req_addr,
  input  [2:0]   io_in_bits_req_size,
  input  [86:0]  io_in_bits_req_user,
  input  [3:0]   io_in_bits_hitVec,
  input          io_in_bits_miss,
  input          io_in_bits_hitWB,
  input          io_in_bits_hitinstrPF,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [86:0]  io_out_bits_user,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input          io_flush,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output         io_ipf,
  output         io_isFinish
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  missIPF; // @[EmbeddedTLB.scala 686:24]
  wire [8:0] vpn_vpn0 = io_in_bits_req_addr[20:12]; // @[EmbeddedTLB.scala 694:54]
  wire [8:0] vpn_vpn1 = io_in_bits_req_addr[29:21]; // @[EmbeddedTLB.scala 694:54]
  wire [8:0] vpn_vpn2 = io_in_bits_req_addr[38:30]; // @[EmbeddedTLB.scala 694:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 696:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 696:30]
  wire  hit = io_in_valid & |io_in_bits_hitVec; // @[EmbeddedTLB.scala 701:25]
  wire  miss = io_in_valid & io_in_bits_miss; // @[EmbeddedTLB.scala 702:26]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_16 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_19 = {_T_16,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[EmbeddedTLB.scala 704:42]
  wire [3:0] waymask = hit ? io_in_bits_hitVec : victimWaymask; // @[EmbeddedTLB.scala 705:20]
  wire  hitinstrPF = io_in_bits_hitinstrPF & io_in_valid; // @[EmbeddedTLB.scala 709:42]
  wire  hitWB = io_in_bits_hitWB & io_in_valid; // @[EmbeddedTLB.scala 710:32]
  wire [120:0] _T_32 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_33 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_34 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_35 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_36 = _T_32 | _T_33; // @[Mux.scala 27:72]
  wire [120:0] _T_37 = _T_36 | _T_34; // @[Mux.scala 27:72]
  wire [120:0] _T_38 = _T_37 | _T_35; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_38[59:52]; // @[EmbeddedTLB.scala 718:70]
  wire [17:0] hitMeta_mask = _T_38[77:60]; // @[EmbeddedTLB.scala 718:70]
  wire [15:0] hitMeta_asid = _T_38[93:78]; // @[EmbeddedTLB.scala 718:70]
  wire [31:0] hitData_pteaddr = _T_38[31:0]; // @[EmbeddedTLB.scala 719:70]
  wire [19:0] hitData_ppn = _T_38[51:32]; // @[EmbeddedTLB.scala 719:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 720:38]
  wire [7:0] _T_70 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 723:79]
  wire [7:0] hitRefillFlag = 8'h40 | _T_70; // @[EmbeddedTLB.scala 723:69]
  wire [39:0] _T_71 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 30:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  reg [2:0] state; // @[EmbeddedTLB.scala 733:22]
  reg [1:0] level; // @[EmbeddedTLB.scala 734:22]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 736:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 738:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 741:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 741:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 742:18]
  wire  _T_83 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  needFlush; // @[EmbeddedTLB.scala 746:26]
  wire  isFlush = needFlush | io_flush; // @[EmbeddedTLB.scala 748:27]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[EmbeddedTLB.scala 746:26 749:{40,52}]
  wire  _GEN_4 = _T_83 & needFlush ? 1'h0 : _GEN_3; // @[EmbeddedTLB.scala 750:{37,49}]
  wire  _T_89 = ~isFlush; // @[EmbeddedTLB.scala 755:13]
  wire [31:0] _T_94 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 30:58]
  wire  _T_96 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_13 = _T_96 ? 3'h2 : state; // @[EmbeddedTLB.scala 733:22 773:{38,46}]
  wire  _GEN_15 = io_flush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 767:22 769:19]
  wire  _GEN_16 = io_flush ? 1'h0 : missIPF; // @[EmbeddedTLB.scala 767:22 770:17 686:24]
  wire [7:0] _T_98 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,
    memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 777:44]
  wire  _T_107 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_110 = level == 2'h3; // @[EmbeddedTLB.scala 785:58]
  wire  _T_111 = level == 2'h2; // @[EmbeddedTLB.scala 785:73]
  wire [8:0] _T_141 = _T_110 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 801:50]
  wire [31:0] _T_143 = {memRdata_ppn,_T_141,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_19 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? 3'h4 : 3'h1; // @[EmbeddedTLB.scala 786:60 787:43 800:19]
  wire  _GEN_20 = ~_T_98[0] | ~_T_98[1] & _T_98[2] | missIPF; // @[EmbeddedTLB.scala 686:24 786:60 788:45]
  wire [31:0] _GEN_21 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? raddr : _T_143; // @[EmbeddedTLB.scala 742:18 786:60 801:19]
  wire  _T_156 = _T_98[0] & ~(io_pf_priviledgeMode == 2'h0 & ~_T_98[4]) & ~(io_pf_priviledgeMode == 2'h1 & _T_98[4]); // @[EmbeddedTLB.scala 804:87]
  wire  _T_157 = _T_156 & _T_98[3]; // @[EmbeddedTLB.scala 805:36]
  wire  _T_162 = ~_T_98[6]; // @[EmbeddedTLB.scala 808:26]
  wire [7:0] _T_171 = {_T_98[7],_T_98[6],_T_98[5],_T_98[4],_T_98[3],_T_98[2],_T_98[1],_T_98[0]}; // @[EmbeddedTLB.scala 810:79]
  wire [7:0] _T_172 = 8'h40 | _T_171; // @[EmbeddedTLB.scala 810:68]
  wire [63:0] _T_173 = io_mem_resp_bits_rdata | 64'h40; // @[EmbeddedTLB.scala 811:50]
  wire  _GEN_22 = ~_T_157 | _T_162 | missIPF; // @[EmbeddedTLB.scala 813:42 814:23 686:24]
  wire  _GEN_24 = ~_T_157 | _T_162 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 813:42 817:30]
  wire [17:0] _T_178 = _T_111 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 832:59]
  wire [17:0] _T_179 = _T_110 ? 18'h0 : _T_178; // @[EmbeddedTLB.scala 832:26]
  wire [7:0] _GEN_25 = level != 2'h0 ? _T_172 : 8'h0; // @[EmbeddedTLB.scala 803:36 810:26]
  wire [63:0] _GEN_26 = level != 2'h0 ? _T_173 : memRespStore; // @[EmbeddedTLB.scala 803:36 811:24 736:25]
  wire  _GEN_27 = level != 2'h0 ? _GEN_22 : missIPF; // @[EmbeddedTLB.scala 686:24 803:36]
  wire [2:0] _GEN_28 = level != 2'h0 ? 3'h4 : state; // @[EmbeddedTLB.scala 733:22 803:36]
  wire  _GEN_29 = level != 2'h0 & _GEN_24; // @[EmbeddedTLB.scala 803:36]
  wire [17:0] _GEN_30 = level != 2'h0 ? _T_179 : 18'h3ffff; // @[EmbeddedTLB.scala 803:36 832:20]
  wire [17:0] _GEN_38 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_30; // @[EmbeddedTLB.scala 785:82]
  wire [17:0] _GEN_49 = isFlush ? 18'h3ffff : _GEN_38; // @[EmbeddedTLB.scala 779:24]
  wire [17:0] _GEN_60 = _T_107 ? _GEN_49 : 18'h3ffff; // @[EmbeddedTLB.scala 778:33]
  wire [17:0] _GEN_111 = 3'h2 == state ? _GEN_60 : 18'h3ffff; // @[EmbeddedTLB.scala 753:18]
  wire [17:0] _GEN_123 = 3'h1 == state ? 18'h3ffff : _GEN_111; // @[EmbeddedTLB.scala 753:18]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_123; // @[EmbeddedTLB.scala 753:18]
  wire [17:0] _GEN_31 = level != 2'h0 ? missMask : missMaskStore; // @[EmbeddedTLB.scala 803:36 833:25 738:26]
  wire [2:0] _GEN_32 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_28; // @[EmbeddedTLB.scala 785:82]
  wire  _GEN_33 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : _GEN_27; // @[EmbeddedTLB.scala 785:82]
  wire [31:0] _GEN_34 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_21 : raddr; // @[EmbeddedTLB.scala 742:18 785:82]
  wire [7:0] _GEN_35 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_25; // @[EmbeddedTLB.scala 785:82]
  wire [63:0] _GEN_36 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_26; // @[EmbeddedTLB.scala 736:25 785:82]
  wire  _GEN_37 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_29; // @[EmbeddedTLB.scala 785:82]
  wire [17:0] _GEN_39 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_31; // @[EmbeddedTLB.scala 738:26 785:82]
  wire [2:0] _GEN_40 = isFlush ? 3'h0 : _GEN_32; // @[EmbeddedTLB.scala 779:24 780:17]
  wire  _GEN_41 = isFlush ? 1'h0 : _GEN_33; // @[EmbeddedTLB.scala 779:24 781:19]
  wire  _GEN_44 = isFlush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 779:24 784:21]
  wire [31:0] _GEN_45 = isFlush ? raddr : _GEN_34; // @[EmbeddedTLB.scala 742:18 779:24]
  wire [7:0] _GEN_46 = isFlush ? 8'h0 : _GEN_35; // @[EmbeddedTLB.scala 779:24]
  wire [63:0] _GEN_47 = isFlush ? memRespStore : _GEN_36; // @[EmbeddedTLB.scala 779:24 736:25]
  wire  _GEN_48 = isFlush ? 1'h0 : _GEN_37; // @[EmbeddedTLB.scala 779:24]
  wire [17:0] _GEN_50 = isFlush ? missMaskStore : _GEN_39; // @[EmbeddedTLB.scala 779:24 738:26]
  wire [1:0] _T_181 = level - 2'h1; // @[EmbeddedTLB.scala 835:24]
  wire [2:0] _GEN_51 = _T_107 ? _GEN_40 : state; // @[EmbeddedTLB.scala 733:22 778:33]
  wire  _GEN_52 = _T_107 ? _GEN_41 : missIPF; // @[EmbeddedTLB.scala 686:24 778:33]
  wire  _GEN_55 = _T_107 ? _GEN_44 : _GEN_4; // @[EmbeddedTLB.scala 778:33]
  wire [7:0] _GEN_57 = _T_107 ? _GEN_46 : 8'h0; // @[EmbeddedTLB.scala 778:33]
  wire  _GEN_59 = _T_107 & _GEN_48; // @[EmbeddedTLB.scala 778:33]
  wire [1:0] _GEN_62 = _T_107 ? _T_181 : level; // @[EmbeddedTLB.scala 778:33 835:15 734:22]
  wire [2:0] _GEN_63 = _T_96 ? 3'h6 : state; // @[EmbeddedTLB.scala 733:22 846:{38,46}]
  wire [2:0] _GEN_64 = io_flush ? 3'h0 : _GEN_63; // @[EmbeddedTLB.scala 840:22 841:15]
  wire [2:0] _GEN_65 = isFlush ? 3'h0 : 3'h4; // @[EmbeddedTLB.scala 851:22 852:17 858:17]
  wire  _GEN_66 = isFlush ? 1'h0 : missIPF; // @[EmbeddedTLB.scala 851:22 854:19 686:24]
  wire [2:0] _GEN_67 = _T_107 ? _GEN_65 : state; // @[EmbeddedTLB.scala 733:22 850:32]
  wire  _GEN_69 = _T_107 ? _GEN_66 : missIPF; // @[EmbeddedTLB.scala 686:24 850:32]
  wire [2:0] _GEN_72 = _T_83 | io_flush ? 3'h0 : state; // @[EmbeddedTLB.scala 863:56 864:13 733:22]
  wire  _GEN_73 = _T_83 | io_flush ? 1'h0 : missIPF; // @[EmbeddedTLB.scala 863:56 865:15 686:24]
  wire  _GEN_76 = _T_83 | io_flush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 863:56 868:17]
  wire [2:0] _GEN_82 = 3'h5 == state ? _GEN_72 : state; // @[EmbeddedTLB.scala 753:18 733:22]
  wire  _GEN_85 = 3'h5 == state ? _GEN_73 : missIPF; // @[EmbeddedTLB.scala 753:18 686:24]
  wire  _GEN_86 = 3'h5 == state ? _GEN_76 : _GEN_4; // @[EmbeddedTLB.scala 753:18]
  wire [2:0] _GEN_87 = 3'h4 == state ? _GEN_72 : _GEN_82; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_88 = 3'h4 == state ? _GEN_73 : _GEN_85; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_91 = 3'h4 == state ? _GEN_76 : _GEN_86; // @[EmbeddedTLB.scala 753:18]
  wire [2:0] _GEN_92 = 3'h6 == state ? _GEN_67 : _GEN_87; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_93 = 3'h6 == state ? _GEN_55 : _GEN_91; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_94 = 3'h6 == state ? _GEN_69 : _GEN_88; // @[EmbeddedTLB.scala 753:18]
  wire [2:0] _GEN_97 = 3'h3 == state ? _GEN_64 : _GEN_92; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_98 = 3'h3 == state ? _GEN_15 : _GEN_93; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_99 = 3'h3 == state ? _GEN_16 : _GEN_94; // @[EmbeddedTLB.scala 753:18]
  wire [7:0] _GEN_108 = 3'h2 == state ? _GEN_57 : 8'h0; // @[EmbeddedTLB.scala 753:18]
  wire [7:0] _GEN_120 = 3'h1 == state ? 8'h0 : _GEN_108; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_122 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_59; // @[EmbeddedTLB.scala 753:18]
  wire [7:0] missRefillFlag = 3'h0 == state ? 8'h0 : _GEN_120; // @[EmbeddedTLB.scala 753:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_122; // @[EmbeddedTLB.scala 753:18]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 883:23]
  wire [31:0] _T_193 = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 884:35]
  wire  _T_198 = ~io_flush; // @[EmbeddedTLB.scala 885:77]
  wire [15:0] _T_212 = hitWB ? hitMeta_asid : satp_asid; // @[EmbeddedTLB.scala 891:15]
  wire [17:0] _T_213 = hitWB ? hitMeta_mask : missMask; // @[EmbeddedTLB.scala 891:59]
  wire [7:0] _T_214 = hitWB ? hitRefillFlag : missRefillFlag; // @[EmbeddedTLB.scala 892:15]
  wire [19:0] _T_215 = hitWB ? hitData_ppn : memRdata_ppn; // @[EmbeddedTLB.scala 892:64]
  wire [59:0] lo_5 = {_T_214,_T_215,_T_193}; // @[Cat.scala 30:58]
  wire [60:0] hi_8 = {vpn_vpn2,vpn_vpn1,vpn_vpn0,_T_212,_T_213}; // @[Cat.scala 30:58]
  wire [31:0] _T_219 = {hitData_ppn,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_221 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_222 = _T_219 & _T_221; // @[BitUtils.scala 32:13]
  wire [31:0] _T_223 = ~_T_221; // @[BitUtils.scala 32:38]
  wire [31:0] _T_224 = io_in_bits_req_addr[31:0] & _T_223; // @[BitUtils.scala 32:36]
  wire [31:0] _T_225 = _T_222 | _T_224; // @[BitUtils.scala 32:25]
  wire [31:0] _T_238 = {memRespStore[29:10],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_240 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_241 = _T_238 & _T_240; // @[BitUtils.scala 32:13]
  wire [31:0] _T_242 = ~_T_240; // @[BitUtils.scala 32:38]
  wire [31:0] _T_243 = io_in_bits_req_addr[31:0] & _T_242; // @[BitUtils.scala 32:36]
  wire [31:0] _T_244 = _T_241 | _T_243; // @[BitUtils.scala 32:25]
  wire  _T_248 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 176:23]
  assign io_in_ready = ~io_in_valid | _T_83 & io_mdReady; // @[EmbeddedTLB.scala 900:31]
  assign io_out_valid = _T_198 & io_in_valid & (state == 3'h4 & ~(_T_248 | io_ipf)); // @[EmbeddedTLB.scala 898:43]
  assign io_out_bits_addr = hit ? _T_225 : _T_244; // @[EmbeddedTLB.scala 897:26]
  assign io_out_bits_size = io_in_bits_req_size; // @[EmbeddedTLB.scala 896:15]
  assign io_out_bits_user = io_in_bits_req_user; // @[EmbeddedTLB.scala 896:15]
  assign io_mdWrite_wen = io_in_valid & (missMetaRefill & _T_89 | hitWB & state == 3'h0 & _T_89); // @[EmbeddedTLB.scala 889:38]
  assign io_mdWrite_waymask = hit ? io_in_bits_hitVec : victimWaymask; // @[EmbeddedTLB.scala 705:20]
  assign io_mdWrite_wdata = {hi_8,lo_5}; // @[Cat.scala 30:58]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~io_flush; // @[EmbeddedTLB.scala 885:74]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 884:35]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[EmbeddedTLB.scala 884:138]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 886:21]
  assign io_pf_loadPF = 1'h0; // @[EmbeddedTLB.scala 713:39]
  assign io_pf_storePF = 1'h0; // @[EmbeddedTLB.scala 714:41]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[EmbeddedTLB.scala 902:16]
  assign io_isFinish = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  always @(posedge clock) begin
    if (reset) begin // @[EmbeddedTLB.scala 686:24]
      missIPF <= 1'h0; // @[EmbeddedTLB.scala 686:24]
    end else if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
        if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
          missIPF <= 1'h0; // @[EmbeddedTLB.scala 770:17]
        end
      end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        missIPF <= _GEN_52;
      end else begin
        missIPF <= _GEN_99;
      end
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_19;
    end
    if (hitWB) begin // @[Reg.scala 16:19]
      hitWBStore <= _T_71; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 733:22]
      state <= 3'h0; // @[EmbeddedTLB.scala 733:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (~isFlush & hitWB) begin // @[EmbeddedTLB.scala 755:32]
        state <= 3'h3; // @[EmbeddedTLB.scala 756:15]
      end else if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
        state <= 3'h1; // @[EmbeddedTLB.scala 759:15]
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
        state <= 3'h0; // @[EmbeddedTLB.scala 768:15]
      end else begin
        state <= _GEN_13;
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
      state <= _GEN_51;
    end else begin
      state <= _GEN_97;
    end
    if (reset) begin // @[EmbeddedTLB.scala 734:22]
      level <= 2'h3; // @[EmbeddedTLB.scala 734:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (!(~isFlush & hitWB)) begin // @[EmbeddedTLB.scala 755:32]
        if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
          level <= 2'h3; // @[EmbeddedTLB.scala 761:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        level <= _GEN_62;
      end
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
          if (_T_107) begin // @[EmbeddedTLB.scala 778:33]
            memRespStore <= _GEN_47;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
          if (_T_107) begin // @[EmbeddedTLB.scala 778:33]
            missMaskStore <= _GEN_50;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (!(~isFlush & hitWB)) begin // @[EmbeddedTLB.scala 755:32]
        if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
          raddr <= _T_94; // @[EmbeddedTLB.scala 760:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        if (_T_107) begin // @[EmbeddedTLB.scala 778:33]
          raddr <= _GEN_45;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 746:26]
      needFlush <= 1'h0; // @[EmbeddedTLB.scala 746:26]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (~isFlush & hitWB) begin // @[EmbeddedTLB.scala 755:32]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 757:19]
      end else if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 762:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 769:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
      needFlush <= _GEN_55;
    end else begin
      needFlush <= _GEN_98;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  missIPF = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  hitWBStore = _RAND_2[39:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  level = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  memRespStore = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  missMaskStore = _RAND_6[17:0];
  _RAND_7 = {1{`RANDOM}};
  raddr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_1 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_2 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_3 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg  resetState; // @[EmbeddedTLB.scala 55:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[EmbeddedTLB.scala 57:22 55:27 57:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 66:20]
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = 1'h0;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = 1'h0;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = 1'h0;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = 1'h0;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = 1'h0;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = 1'h0;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = 1'h0;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = 1'h0;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 72:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    resetState <= reset | _GEN_1; // @[EmbeddedTLB.scala 55:{27,27}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SIMD_TLB(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [86:0] io_out_req_bits_user,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input  [86:0] io_out_resp_bits_user,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_flush,
  input  [1:0]  io_csrMMU_priviledgeMode,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  input         io_cacheEmpty,
  output        io_ipf,
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 443:23]
  wire [38:0] tlbExec_io_in_bits_req_addr; // @[EmbeddedTLB.scala 443:23]
  wire [2:0] tlbExec_io_in_bits_req_size; // @[EmbeddedTLB.scala 443:23]
  wire [86:0] tlbExec_io_in_bits_req_user; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_in_bits_hitVec; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_miss; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_hitWB; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_hitinstrPF; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 443:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 443:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 443:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 443:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_flush; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 443:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 443:23]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 445:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 445:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 445:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 445:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 445:21]
  reg [120:0] r__0; // @[Reg.scala 15:16]
  reg [120:0] r__1; // @[Reg.scala 15:16]
  reg [120:0] r__2; // @[Reg.scala 15:16]
  reg [120:0] r__3; // @[Reg.scala 15:16]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 470:57]
  wire [120:0] _WIRE_46 = mdTLB_io_tlbmd_3;
  wire [26:0] _T_205 = {9'h1ff,_WIRE_46[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_206 = _T_205 & _WIRE_46[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_204 = {io_in_req_bits_addr[38:30],io_in_req_bits_addr[29:21],io_in_req_bits_addr[20:12]}; // @[EmbeddedTLB.scala 531:224]
  wire [26:0] _T_208 = _T_205 & _T_204; // @[TLB.scala 131:84]
  wire  _T_209 = _T_206 == _T_208; // @[TLB.scala 131:48]
  wire  _T_210 = _WIRE_46[52] & _WIRE_46[93:78] == CSRSATP[59:44] & _T_209; // @[EmbeddedTLB.scala 531:155]
  wire [120:0] _WIRE_34 = mdTLB_io_tlbmd_2;
  wire [26:0] _T_160 = {9'h1ff,_WIRE_34[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_161 = _T_160 & _WIRE_34[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_163 = _T_160 & _T_204; // @[TLB.scala 131:84]
  wire  _T_164 = _T_161 == _T_163; // @[TLB.scala 131:48]
  wire  _T_165 = _WIRE_34[52] & _WIRE_34[93:78] == CSRSATP[59:44] & _T_164; // @[EmbeddedTLB.scala 531:155]
  wire [120:0] _WIRE_22 = mdTLB_io_tlbmd_1;
  wire [26:0] _T_115 = {9'h1ff,_WIRE_22[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_116 = _T_115 & _WIRE_22[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_118 = _T_115 & _T_204; // @[TLB.scala 131:84]
  wire  _T_119 = _T_116 == _T_118; // @[TLB.scala 131:48]
  wire  _T_120 = _WIRE_22[52] & _WIRE_22[93:78] == CSRSATP[59:44] & _T_119; // @[EmbeddedTLB.scala 531:155]
  wire [120:0] _WIRE_10 = mdTLB_io_tlbmd_0;
  wire [26:0] _T_70 = {9'h1ff,_WIRE_10[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_71 = _T_70 & _WIRE_10[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_73 = _T_70 & _T_204; // @[TLB.scala 131:84]
  wire  _T_74 = _T_71 == _T_73; // @[TLB.scala 131:48]
  wire  _T_75 = _WIRE_10[52] & _WIRE_10[93:78] == CSRSATP[59:44] & _T_74; // @[EmbeddedTLB.scala 531:155]
  wire [3:0] _T_211 = {_T_210,_T_165,_T_120,_T_75}; // @[EmbeddedTLB.scala 531:234]
  wire  _T_214 = |_T_211; // @[EmbeddedTLB.scala 533:43]
  wire  _T_216 = io_in_req_valid & ~(|_T_211); // @[EmbeddedTLB.scala 533:32]
  wire  _T_213 = io_in_req_valid & _T_214; // @[EmbeddedTLB.scala 532:31]
  reg [63:0] REG_4; // @[LFSR64.scala 25:23]
  wire [3:0] _T_229 = 4'h1 << REG_4[1:0]; // @[EmbeddedTLB.scala 535:44]
  wire [3:0] _T_230 = _T_213 ? _T_211 : _T_229; // @[EmbeddedTLB.scala 536:22]
  wire [120:0] _T_235 = _T_230[0] ? mdTLB_io_tlbmd_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_236 = _T_230[1] ? mdTLB_io_tlbmd_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_239 = _T_235 | _T_236; // @[Mux.scala 27:72]
  wire [120:0] _T_237 = _T_230[2] ? mdTLB_io_tlbmd_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_240 = _T_239 | _T_237; // @[Mux.scala 27:72]
  wire [120:0] _T_238 = _T_230[3] ? mdTLB_io_tlbmd_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_241 = _T_240 | _T_238; // @[Mux.scala 27:72]
  wire  _T_300 = _T_213 & ~(io_csrMMU_priviledgeMode == 2'h0 & ~_T_241[56]) & ~(io_csrMMU_priviledgeMode == 2'h1 &
    _T_241[56]); // @[EmbeddedTLB.scala 557:96]
  wire  _T_301 = _T_300 & _T_241[55]; // @[EmbeddedTLB.scala 558:28]
  wire  _T_307 = ~_T_301 & _T_213; // @[EmbeddedTLB.scala 570:54]
  wire  _T_280 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 176:23]
  wire  _T_282 = ~_T_280; // @[EmbeddedTLB.scala 552:86]
  wire  _T_283 = _T_213 & ~_T_241[58] & ~_T_307 & ~_T_280; // @[EmbeddedTLB.scala 552:83]
  wire  _T_350 = _T_216 | _T_283 | _T_307; // @[EmbeddedTLB.scala 609:86]
  wire  tlbexec_inbundle_valid = ~vmEnable ? 1'h0 : io_in_req_valid & (_T_216 | _T_283 | _T_307); // @[EmbeddedTLB.scala 507:19 508:28 609:28]
  wire  mdUpdate = tlbexec_inbundle_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 482:26]
  reg  REG_3; // @[EmbeddedTLB.scala 473:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : REG_3; // @[EmbeddedTLB.scala 473:24 474:{25,33}]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[EmbeddedTLB.scala 475:{50,58}]
  reg [38:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_1_req_size; // @[Reg.scala 15:16]
  reg [86:0] r_1_req_user; // @[Reg.scala 15:16]
  reg [3:0] r_1_hitVec; // @[Reg.scala 15:16]
  reg  r_1_miss; // @[Reg.scala 15:16]
  reg  r_1_hitWB; // @[Reg.scala 15:16]
  reg  r_1_hitinstrPF; // @[Reg.scala 15:16]
  reg  state; // @[EmbeddedTLB.scala 505:22]
  wire  _T_223 = REG_4[0] ^ REG_4[1] ^ REG_4[3] ^ REG_4[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_226 = {_T_223,REG_4[63:1]}; // @[Cat.scala 30:58]
  wire  _T_308 = ~state; // @[EmbeddedTLB.scala 577:32]
  wire  _T_316 = ~state ? _T_213 & ~_T_283 & _T_282 : tlbExec_io_out_valid; // @[EmbeddedTLB.scala 577:25]
  wire [31:0] _T_319 = {_T_241[51:32],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_321 = {2'h3,_T_241[77:60],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_322 = _T_319 & _T_321; // @[BitUtils.scala 32:13]
  wire [31:0] _T_323 = ~_T_321; // @[BitUtils.scala 32:38]
  wire [31:0] _T_324 = io_in_req_bits_addr[31:0] & _T_323; // @[BitUtils.scala 32:36]
  wire [31:0] _T_325 = _T_322 | _T_324; // @[BitUtils.scala 32:25]
  wire [31:0] _T_326 = _T_308 ? _T_325 : tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 578:29]
  wire  out_req_ready = ~vmEnable ? 1'h0 : io_out_req_ready; // @[EmbeddedTLB.scala 507:19 522:19 583:19]
  wire  _T_376 = tlbExec_io_ipf & vmEnable; // @[EmbeddedTLB.scala 639:26]
  wire  _GEN_43 = ~vmEnable ? 1'h0 : _T_316; // @[EmbeddedTLB.scala 507:19 521:19 577:19]
  wire  out_req_valid = tlbExec_io_ipf & vmEnable ? 1'h0 : _GEN_43; // @[EmbeddedTLB.scala 639:39 641:21]
  wire  _T_327 = out_req_ready & out_req_valid; // @[Decoupled.scala 40:37]
  wire  tlbexec_inbundle_ready = tlbExec_io_in_ready; // @[EmbeddedTLB.scala 478:16 490:30]
  wire  _T_336 = tlbexec_inbundle_ready & tlbexec_inbundle_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_22 = _T_350 & ~io_flush & _T_336 | state; // @[EmbeddedTLB.scala 588:105 589:17 505:22]
  wire  _GEN_23 = _T_327 | io_flush ? 1'h0 : state; // @[EmbeddedTLB.scala 593:41 595:17 505:22]
  wire  _GEN_24 = ~io_in_req_valid ? 1'h0 : _GEN_23; // @[EmbeddedTLB.scala 597:31 598:17]
  wire  _GEN_25 = ~io_in_req_valid | io_flush; // @[EmbeddedTLB.scala 448:20 597:31 599:28]
  wire  _GEN_27 = state ? _GEN_25 : io_flush; // @[EmbeddedTLB.scala 586:19 448:20]
  wire  _GEN_29 = _T_308 ? io_flush : _GEN_27; // @[EmbeddedTLB.scala 586:19 448:20]
  wire [31:0] _GEN_51 = ~vmEnable ? tlbExec_io_out_bits_addr : _T_326; // @[EmbeddedTLB.scala 495:16 507:19 578:23]
  wire [38:0] out_req_bits_addr = {{7'd0}, _GEN_51}; // @[EmbeddedTLB.scala 494:21]
  wire  _GEN_33 = ~vmEnable | _T_327; // @[EmbeddedTLB.scala 507:19 509:26 579:26]
  wire [38:0] _GEN_36 = ~vmEnable ? {{7'd0}, io_in_req_bits_addr[31:0]} : out_req_bits_addr; // @[EmbeddedTLB.scala 507:19 514:26 583:19]
  wire [2:0] out_req_bits_size = ~vmEnable ? tlbExec_io_out_bits_size : 3'h3; // @[EmbeddedTLB.scala 495:16 507:19 576:18]
  wire [86:0] out_req_bits_user = ~vmEnable ? tlbExec_io_out_bits_user : io_in_req_bits_user; // @[EmbeddedTLB.scala 495:16 507:19 576:18]
  SIMD_TLBEXEC tlbExec ( // @[EmbeddedTLB.scala 443:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_req_addr(tlbExec_io_in_bits_req_addr),
    .io_in_bits_req_size(tlbExec_io_in_bits_req_size),
    .io_in_bits_req_user(tlbExec_io_in_bits_req_user),
    .io_in_bits_hitVec(tlbExec_io_in_bits_hitVec),
    .io_in_bits_miss(tlbExec_io_in_bits_miss),
    .io_in_bits_hitWB(tlbExec_io_in_bits_hitWB),
    .io_in_bits_hitinstrPF(tlbExec_io_in_bits_hitinstrPF),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  EmbeddedTLBMD mdTLB ( // @[EmbeddedTLB.scala 445:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : _T_327; // @[EmbeddedTLB.scala 507:19 513:21 580:21]
  assign io_in_resp_valid = _T_376 & io_cacheEmpty | io_out_resp_valid; // @[EmbeddedTLB.scala 620:14 644:56 645:24]
  assign io_in_resp_bits_rdata = _T_376 & io_cacheEmpty ? 64'h0 : io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 620:14 644:56 646:29]
  assign io_in_resp_bits_user = _T_376 & io_cacheEmpty ? tlbExec_io_in_bits_req_user : io_out_resp_bits_user; // @[EmbeddedTLB.scala 620:14 644:56 648:34]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : out_req_valid; // @[EmbeddedTLB.scala 507:19 512:22 583:19]
  assign io_out_req_bits_addr = _GEN_36[31:0];
  assign io_out_req_bits_size = ~vmEnable ? 3'h3 : out_req_bits_size; // @[EmbeddedTLB.scala 507:19 515:26 583:19]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : out_req_bits_user; // @[EmbeddedTLB.scala 507:19 519:32 583:19]
  assign io_out_resp_ready = io_in_resp_ready; // @[EmbeddedTLB.scala 620:14]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 450:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 450:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 450:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 450:18]
  assign io_csrMMU_loadPF = 1'h0; // @[EmbeddedTLB.scala 454:20]
  assign io_csrMMU_storePF = 1'h0; // @[EmbeddedTLB.scala 455:21]
  assign io_ipf = _T_376 & io_cacheEmpty & tlbExec_io_ipf; // @[EmbeddedTLB.scala 462:10 644:56 649:14]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = REG_3; // @[EmbeddedTLB.scala 480:17]
  assign tlbExec_io_in_bits_req_addr = r_1_req_addr; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_req_size = r_1_req_size; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_req_user = r_1_req_user; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_hitVec = r_1_hitVec; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_miss = r_1_miss; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_hitWB = r_1_hitWB; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_hitinstrPF = r_1_hitinstrPF; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_out_ready = tlbExec_io_ipf & vmEnable ? io_cacheEmpty & io_in_resp_ready : _GEN_33; // @[EmbeddedTLB.scala 639:39 640:28]
  assign tlbExec_io_md_0 = r__0; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_md_1 = r__1; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_md_2 = r__2; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_md_3 = r__3; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 458:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 450:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 450:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 450:18]
  assign tlbExec_io_flush = ~vmEnable ? io_flush : _GEN_29; // @[EmbeddedTLB.scala 507:19 448:20]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 449:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 451:32]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 467:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 460:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 460:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 460:18]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__0 <= mdTLB_io_tlbmd_0; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__1 <= mdTLB_io_tlbmd_1; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__2 <= mdTLB_io_tlbmd_2; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__3 <= mdTLB_io_tlbmd_3; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG_4 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG_4 == 64'h0) begin // @[LFSR64.scala 28:18]
      REG_4 <= 64'h1;
    end else begin
      REG_4 <= _T_226;
    end
    if (reset) begin // @[EmbeddedTLB.scala 473:24]
      REG_3 <= 1'h0; // @[EmbeddedTLB.scala 473:24]
    end else if (io_flush) begin // @[EmbeddedTLB.scala 476:20]
      REG_3 <= 1'h0; // @[EmbeddedTLB.scala 476:28]
    end else begin
      REG_3 <= _GEN_5;
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_addr <= 39'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_addr <= io_in_req_bits_addr; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_size <= 3'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_size <= 3'h3; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_user <= 87'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_user <= io_in_req_bits_user; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_hitVec <= 4'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_hitVec <= _T_211; // @[EmbeddedTLB.scala 610:34]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_miss <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_miss <= _T_216; // @[EmbeddedTLB.scala 611:32]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_hitWB <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_hitWB <= _T_283; // @[EmbeddedTLB.scala 612:33]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_hitinstrPF <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_hitinstrPF <= _T_307; // @[EmbeddedTLB.scala 615:38]
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 505:22]
      state <= 1'h0; // @[EmbeddedTLB.scala 505:22]
    end else if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
      if (io_flush) begin // @[EmbeddedTLB.scala 520:19]
        state <= 1'h0; // @[EmbeddedTLB.scala 520:26]
      end
    end else if (_T_308) begin // @[EmbeddedTLB.scala 586:19]
      state <= _GEN_22;
    end else if (state) begin // @[EmbeddedTLB.scala 586:19]
      state <= _GEN_24;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  r__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  r__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  r__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  r__3 = _RAND_3[120:0];
  _RAND_4 = {2{`RANDOM}};
  REG_4 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_3 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_req_addr = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_req_size = _RAND_7[2:0];
  _RAND_8 = {3{`RANDOM}};
  r_1_req_user = _RAND_8[86:0];
  _RAND_9 = {1{`RANDOM}};
  r_1_hitVec = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_miss = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_1_hitWB = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_1_hitinstrPF = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [86:0] io_in_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [86:0] io_out_bits_req_user,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_30 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_30) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 147:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 146:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 145:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 145:19]
  assign io_out_bits_req_user = io_in_bits_user; // @[Cache.scala 145:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module CacheStage2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [86:0] io_in_bits_req_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [86:0] io_out_bits_req_user,
  output [18:0] io_out_bits_metas_0_tag,
  output [18:0] io_out_bits_metas_1_tag,
  output [18:0] io_out_bits_metas_2_tag,
  output [18:0] io_out_bits_metas_3_tag,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 176:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 176:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 176:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 178:64]
  reg  isForwardMetaReg; // @[Cache.scala 179:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 180:24 179:33 180:43]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 181:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 181:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 15:16 16:{19,23}]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 15:16 16:{19,23}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 185:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 187:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 187:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 187:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 187:61]
  wire [18:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[Cache.scala 189:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 192:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_39 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_42 = {_T_39,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 193:42]
  wire  _T_45 = ~metaWay_0_valid; // @[Cache.scala 195:45]
  wire  _T_46 = ~metaWay_1_valid; // @[Cache.scala 195:45]
  wire  _T_47 = ~metaWay_2_valid; // @[Cache.scala 195:45]
  wire  _T_48 = ~metaWay_3_valid; // @[Cache.scala 195:45]
  wire [3:0] invalidVec = {_T_48,_T_47,_T_46,_T_45}; // @[Cache.scala 195:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 196:34]
  wire [1:0] _T_52 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 199:8]
  wire [2:0] _T_53 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_52}; // @[Cache.scala 198:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_53}; // @[Cache.scala 197:33]
  wire [3:0] _T_54 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 202:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  wire [1:0] _T_59 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_61 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_63 = _T_59 + _T_61; // @[Bitwise.scala 47:55]
  wire  _T_65 = _T_63 > 3'h1; // @[Cache.scala 203:26]
  wire  _T_173 = io_in_bits_req_addr < 32'h40000000; // @[NutCore.scala 92:35]
  wire  _T_177 = io_in_bits_req_addr >= 32'h40600000 & io_in_bits_req_addr < 32'h41600000; // @[NutCore.scala 92:26]
  wire [9:0] _T_194 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_196 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_194; // @[Cache.scala 220:13]
  wire  isForwardData = io_in_valid & _T_196; // @[Cache.scala 219:35]
  reg  isForwardDataReg; // @[Cache.scala 222:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 223:24 222:33 223:43]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_203 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_203; // @[Cache.scala 231:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 230:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 229:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 229:19]
  assign io_out_bits_req_user = io_in_bits_req_user; // @[Cache.scala 229:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 215:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 213:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  assign io_out_bits_mmio = _T_173 | _T_177; // @[NutCore.scala 93:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 226:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 227:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 227:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 179:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 179:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 181:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 181:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_42;
    end
    if (reset) begin // @[Cache.scala 222:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 222:33]
    end else if (_T_12) begin // @[Cache.scala 224:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 224:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 16:23]
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:210 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 210:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fatal; // @[Cache.scala 210:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  REG = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  isForwardDataReg = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_6[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_setIdx,
  input  [18:0] io_in_0_bits_data_tag,
  input         io_in_0_bits_data_dirty,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [6:0]  io_in_1_bits_setIdx,
  input  [18:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [6:0]  io_out_bits_setIdx,
  output [18:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid ? io_in_0_bits_data_dirty : io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module Arbiter_1(
  input         io_in_0_valid,
  input  [9:0]  io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [9:0]  io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [9:0]  io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module CacheStage3(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [86:0] io_in_bits_req_user,
  input  [18:0] io_in_bits_metas_0_tag,
  input  [18:0] io_in_bits_metas_1_tag,
  input  [18:0] io_in_bits_metas_2_tag,
  input  [18:0] io_in_bits_metas_3_tag,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_rdata,
  output [86:0] io_out_bits_user,
  output        io_isFinish,
  input         io_flush,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 257:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 257:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 257:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 257:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 257:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 257:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 258:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 258:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 258:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 258:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 258:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 258:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 261:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 261:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 262:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 263:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 264:26]
  wire [18:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [18:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 277:49]
  wire [63:0] _T_50 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_51 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_52 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_53 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_54 = _T_50 | _T_51; // @[Mux.scala 27:72]
  wire [63:0] _T_55 = _T_54 | _T_52; // @[Mux.scala 27:72]
  wire [63:0] _T_56 = _T_55 | _T_53; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_56; // @[Cache.scala 279:21]
  wire  _T_85 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [3:0] state; // @[Cache.scala 298:22]
  reg  needFlush; // @[Cache.scala 299:26]
  wire  _GEN_1 = io_flush & state != 4'h0 | needFlush; // @[Cache.scala 299:26 301:{41,53}]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 308:23]
  wire  _T_110 = state == 4'h3; // @[Cache.scala 310:39]
  wire  _T_111 = state == 4'h8; // @[Cache.scala 310:66]
  wire [2:0] _T_116 = _T_111 ? value_1 : value_2; // @[Cache.scala 311:33]
  wire  _T_118 = state2 == 2'h1; // @[Cache.scala 312:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_123 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_124 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_125 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_126 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_127 = _T_123 | _T_124; // @[Mux.scala 27:72]
  wire [63:0] _T_128 = _T_127 | _T_125; // @[Mux.scala 27:72]
  wire  _T_131 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_134 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_8 = _T_134 | io_cohResp_valid ? 2'h0 : state2; // @[Cache.scala 318:{100,109} 308:23]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_140 = state == 4'h1; // @[Cache.scala 326:23]
  wire [2:0] _T_142 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 327:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_142; // @[Cache.scala 326:16]
  wire  _T_148 = state2 == 2'h2; // @[Cache.scala 333:89]
  reg  afterFirstRead; // @[Cache.scala 340:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_85 | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_154 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_156 = state == 4'h2; // @[Cache.scala 342:70]
  wire  readingFirst = ~afterFirstRead & _T_154 & state == 4'h2; // @[Cache.scala 342:60]
  wire  _T_159 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 344:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_160 = state == 4'h0; // @[Cache.scala 347:31]
  wire  _T_194 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_196 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = _T_196 ? 4'h7 : state; // @[Cache.scala 298:22 376:{50,58}]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid ? _value_T_7 : value_1; // @[Cache.scala 379:48 Counter.scala 76:15 60:40]
  wire [3:0] _GEN_29 = _T_134 ? 4'h2 : state; // @[Cache.scala 383:50 384:13 298:22]
  wire [2:0] _GEN_30 = _T_134 ? addr_wordIndex : value_1; // @[Cache.scala 383:50 385:25 Counter.scala 60:40]
  wire  _T_210 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_210 ? 4'h7 : state; // @[Cache.scala 298:22 393:{46,54}]
  wire  _GEN_33 = _T_154 | afterFirstRead; // @[Cache.scala 389:33 390:24 340:31]
  wire [2:0] _GEN_34 = _T_154 ? _value_T_7 : value_1; // @[Cache.scala 389:33 Counter.scala 76:15 60:40]
  wire [3:0] _GEN_36 = _T_154 ? _GEN_32 : state; // @[Cache.scala 298:22 389:33]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_134 ? _value_T_11 : value_2; // @[Cache.scala 398:32 Counter.scala 76:15 60:40]
  wire  _T_213 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_213 & _T_134 ? 4'h4 : state; // @[Cache.scala 298:22 399:{65,73}]
  wire [3:0] _GEN_39 = _T_154 ? 4'h1 : state; // @[Cache.scala 298:22 402:{53,61}]
  wire [3:0] _GEN_40 = _T_85 | needFlush | alreadyOutFire ? 4'h0 : state; // @[Cache.scala 298:22 403:{76,84}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[Cache.scala 357:18 298:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[Cache.scala 357:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : value_2; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[Cache.scala 357:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : value_1; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[Cache.scala 357:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? value_2 : _GEN_43; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[Cache.scala 357:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[Cache.scala 357:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_54 = 4'h1 == state ? value_2 : _GEN_49; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[Cache.scala 357:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? state : _GEN_50; // @[Cache.scala 357:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_59 = 4'h8 == state ? value_2 : _GEN_54; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire  dataRefillWriteBus_req_valid = _T_156 & _T_154; // @[Cache.scala 408:39]
  wire  _T_255 = state == 4'h7; // @[Cache.scala 450:48]
  wire  _T_274 = mmio ? _T_255 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 451:45]
  wire  _T_275 = hit | _T_274; // @[Cache.scala 451:28]
  Arbiter metaWriteArb ( // @[Cache.scala 257:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 258:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & _T_160 & ~miss; // @[Cache.scala 462:70]
  assign io_out_valid = io_in_valid & _T_275; // @[Cache.scala 449:31]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 443:29]
  assign io_out_bits_user = io_in_bits_req_user; // @[Cache.scala 446:56]
  assign io_isFinish = hit ? _T_85 : _T_255 & _GEN_12; // @[Cache.scala 459:8]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 310:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_116}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 413:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 423:23]
  assign io_mem_req_valid = _T_140 | _T_110 & state2 == 2'h2; // @[Cache.scala 333:48]
  assign io_mem_req_bits_addr = _T_140 ? raddr : waddr; // @[Cache.scala 328:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_128 | _T_126; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 332:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 338:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 336:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 336:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 337:22]
  assign io_cohResp_valid = _T_111 & _T_148; // @[Cache.scala 348:46]
  assign metaWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 293:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h0; // @[Cache.scala 294:16 97:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 292:29 SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_210; // @[Cache.scala 416:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 261:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = 1'h0; // @[Cache.scala 417:85]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 415:32 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 287:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = useForwardData ? io_in_bits_forwardData_data_data : _T_56; // @[Cache.scala 279:21]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 288:29 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _T_156 & _T_154; // @[Cache.scala 408:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = io_mem_resp_bits_rdata; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 407:32 SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 298:22]
      state <= 4'h0; // @[Cache.scala 298:22]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      if ((miss | mmio) & ~io_flush) begin // @[Cache.scala 370:49]
        if (mmio) begin // @[Cache.scala 371:21]
          state <= 4'h5;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (4'h5 == state) begin // @[Cache.scala 357:18]
      if (_T_194) begin // @[Cache.scala 375:48]
        state <= 4'h6; // @[Cache.scala 375:56]
      end
    end else if (4'h6 == state) begin // @[Cache.scala 357:18]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[Cache.scala 299:26]
      needFlush <= 1'h0; // @[Cache.scala 299:26]
    end else if (_T_85 & needFlush) begin // @[Cache.scala 302:37]
      needFlush <= 1'h0; // @[Cache.scala 302:49]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
          value_1 <= _GEN_55;
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 308:23]
      state2 <= 2'h0; // @[Cache.scala 308:23]
    end else if (2'h0 == state2) begin // @[Cache.scala 315:19]
      if (_T_131) begin // @[Cache.scala 316:53]
        state2 <= 2'h1; // @[Cache.scala 316:62]
      end
    end else if (2'h1 == state2) begin // @[Cache.scala 315:19]
      state2 <= 2'h2; // @[Cache.scala 317:35]
    end else if (2'h2 == state2) begin // @[Cache.scala 315:19]
      state2 <= _GEN_8;
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Cache.scala 340:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 340:31]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      afterFirstRead <= 1'h0; // @[Cache.scala 359:22]
    end else if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      alreadyOutFire <= 1'h0; // @[Cache.scala 360:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_159) begin // @[Reg.scala 16:19]
      if (mmio) begin // @[Cache.scala 343:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:268 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 268:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 268:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  needFlush = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_1(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [6:0]  io_rreq_bits_setIdx,
  output [18:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [18:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [18:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [18:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [18:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  reg  REG; // @[SRAMTemplate.scala 80:30]
  reg [6:0] value; // @[Counter.scala 60:40]
  wire  wrap_wrap = value == 7'h7f; // @[Counter.scala 72:24]
  wire [6:0] _wrap_value_T_1 = value + 7'h1; // @[Counter.scala 76:24]
  wire  wrap = REG & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = wrap ? 1'h0 : REG; // @[SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  wire  _T = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
  wire [6:0] setIdx = REG ? value : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [20:0] _T_1 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = REG ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [20:0] _WIRE_2 = array_RW0_rdata_0;
  wire [20:0] _WIRE_3 = array_RW0_rdata_1;
  wire [20:0] _WIRE_4 = array_RW0_rdata_2;
  wire [20:0] _WIRE_5 = array_RW0_rdata_3;
  array_0 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~REG & _T; // @[SRAMTemplate.scala 101:33]
  assign io_rresp_data_0_tag = _WIRE_2[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_valid = _WIRE_2[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_dirty = _WIRE_2[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_tag = _WIRE_3[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_valid = _WIRE_3[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_dirty = _WIRE_3[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_tag = _WIRE_4[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_valid = _WIRE_4[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_dirty = _WIRE_4[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_tag = _WIRE_5[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_valid = _WIRE_5[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_dirty = _WIRE_5[0]; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | wen;
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[Counter.scala 60:40]
      value <= 7'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      value <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_2(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [6:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [6:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [6:0]  io_r0_req_bits_setIdx,
  output [18:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [18:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [18:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [18:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [18:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [18:0] r_0_tag; // @[Reg.scala 27:20]
  reg  r_0_valid; // @[Reg.scala 27:20]
  reg  r_0_dirty; // @[Reg.scala 27:20]
  reg [18:0] r_1_tag; // @[Reg.scala 27:20]
  reg  r_1_valid; // @[Reg.scala 27:20]
  reg  r_1_dirty; // @[Reg.scala 27:20]
  reg [18:0] r_2_tag; // @[Reg.scala 27:20]
  reg  r_2_valid; // @[Reg.scala 27:20]
  reg  r_2_dirty; // @[Reg.scala 27:20]
  reg [18:0] r_3_tag; // @[Reg.scala 27:20]
  reg  r_3_valid; // @[Reg.scala 27:20]
  reg  r_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_1 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_2 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_tag = REG ? ram_io_rresp_data_0_tag : r_0_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_valid = REG ? ram_io_rresp_data_0_valid : r_0_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_dirty = REG ? ram_io_rresp_data_0_dirty : r_0_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_tag = REG ? ram_io_rresp_data_1_tag : r_1_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_valid = REG ? ram_io_rresp_data_1_valid : r_1_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_dirty = REG ? ram_io_rresp_data_1_dirty : r_1_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_tag = REG ? ram_io_rresp_data_2_tag : r_2_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_valid = REG ? ram_io_rresp_data_2_valid : r_2_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_dirty = REG ? ram_io_rresp_data_2_dirty : r_2_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_tag = REG ? ram_io_rresp_data_3_tag : r_3_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_valid = REG ? ram_io_rresp_data_3_valid : r_3_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_dirty = REG ? ram_io_rresp_data_3_dirty : r_3_dirty; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_0_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_tag <= ram_io_rresp_data_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_valid <= ram_io_rresp_data_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_dirty <= ram_io_rresp_data_0_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_tag <= ram_io_rresp_data_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_valid <= ram_io_rresp_data_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_dirty <= ram_io_rresp_data_1_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_tag <= ram_io_rresp_data_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_valid <= ram_io_rresp_data_2_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_dirty <= ram_io_rresp_data_2_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_tag <= ram_io_rresp_data_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_valid <= ram_io_rresp_data_3_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_dirty <= ram_io_rresp_data_3_dirty; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_0_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  r_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_tag = _RAND_4[18:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_2_tag = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  r_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_3_tag = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  r_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_2(
  input         clock,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [9:0]  io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [9:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire [9:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  wire  realRen = io_rreq_valid & ~io_wreq_valid; // @[SRAMTemplate.scala 89:38]
  array_1 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 101:53]
  assign io_rresp_data_0_data = array_RW0_rdata_0; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_data = array_RW0_rdata_1; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_data = array_RW0_rdata_2; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_data = array_RW0_rdata_3; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = io_wreq_bits_waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = io_wreq_bits_waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = io_wreq_bits_waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = io_wreq_bits_waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | io_wreq_valid;
  assign array_RW0_wmode = io_wreq_valid; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx;
endmodule
module Arbiter_3(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [9:0] io_in_0_bits_setIdx,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [9:0] io_in_1_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [9:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module SRAMTemplateWithArbiter_1(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [9:0]  io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [9:0]  io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [9:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r__0_data; // @[Reg.scala 27:20]
  reg [63:0] r__1_data; // @[Reg.scala 27:20]
  reg [63:0] r__2_data; // @[Reg.scala 27:20]
  reg [63:0] r__3_data; // @[Reg.scala 27:20]
  reg  REG_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r_1_0_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_1_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_2_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_2 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_3 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_data = REG ? ram_io_rresp_data_0_data : r__0_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_data = REG ? ram_io_rresp_data_1_data : r__1_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_data = REG ? ram_io_rresp_data_2_data : r__2_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_data = REG ? ram_io_rresp_data_3_data : r__3_data; // @[Hold.scala 23:48]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r1_resp_data_0_data = REG_1 ? ram_io_rresp_data_0_data : r_1_0_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_1_data = REG_1 ? ram_io_rresp_data_1_data : r_1_1_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_2_data = REG_1 ? ram_io_rresp_data_2_data : r_1_2_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_3_data = REG_1 ? ram_io_rresp_data_3_data : r_1_3_data; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r__0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
    REG_1 <= io_r1_req_ready & io_r1_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_1_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r__0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r__1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  r__2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  r__3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  r_1_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  r_1_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_4(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [86:0] io_in_0_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [86:0] io_out_bits_user
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
  assign io_out_bits_size = io_in_0_bits_size; // @[Arbiter.scala 124:15]
  assign io_out_bits_user = io_in_0_bits_user; // @[Arbiter.scala 124:15]
endmodule
module Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input  [1:0]  io_flush,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_empty,
  input         MOUFlushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 484:18]
  wire  s1_io_in_valid; // @[Cache.scala 484:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 484:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 484:18]
  wire [86:0] s1_io_in_bits_user; // @[Cache.scala 484:18]
  wire  s1_io_out_ready; // @[Cache.scala 484:18]
  wire  s1_io_out_valid; // @[Cache.scala 484:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 484:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 484:18]
  wire [86:0] s1_io_out_bits_req_user; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 484:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 484:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 484:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 484:18]
  wire  s2_clock; // @[Cache.scala 485:18]
  wire  s2_reset; // @[Cache.scala 485:18]
  wire  s2_io_in_ready; // @[Cache.scala 485:18]
  wire  s2_io_in_valid; // @[Cache.scala 485:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 485:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 485:18]
  wire [86:0] s2_io_in_bits_req_user; // @[Cache.scala 485:18]
  wire  s2_io_out_ready; // @[Cache.scala 485:18]
  wire  s2_io_out_valid; // @[Cache.scala 485:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 485:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 485:18]
  wire [86:0] s2_io_out_bits_req_user; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 485:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 485:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 485:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 485:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 485:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 485:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 485:18]
  wire  s3_clock; // @[Cache.scala 486:18]
  wire  s3_reset; // @[Cache.scala 486:18]
  wire  s3_io_in_ready; // @[Cache.scala 486:18]
  wire  s3_io_in_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 486:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 486:18]
  wire [86:0] s3_io_in_bits_req_user; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 486:18]
  wire  s3_io_out_ready; // @[Cache.scala 486:18]
  wire  s3_io_out_valid; // @[Cache.scala 486:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 486:18]
  wire [86:0] s3_io_out_bits_user; // @[Cache.scala 486:18]
  wire  s3_io_isFinish; // @[Cache.scala 486:18]
  wire  s3_io_flush; // @[Cache.scala 486:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 486:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 486:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 486:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 486:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 486:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 486:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 486:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 486:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 486:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 486:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 486:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 486:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 486:18]
  wire  metaArray_clock; // @[Cache.scala 487:25]
  wire  metaArray_reset; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 487:25]
  wire [6:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 487:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 487:25]
  wire [6:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 487:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 487:25]
  wire  dataArray_clock; // @[Cache.scala 488:25]
  wire  dataArray_reset; // @[Cache.scala 488:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 488:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 488:25]
  wire [9:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 488:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 488:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 488:25]
  wire [9:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 488:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 488:25]
  wire [9:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 488:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 488:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 497:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 497:19]
  wire [86:0] arb_io_in_0_bits_user; // @[Cache.scala 497:19]
  wire  arb_io_out_ready; // @[Cache.scala 497:19]
  wire  arb_io_out_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 497:19]
  wire [86:0] arb_io_out_bits_user; // @[Cache.scala 497:19]
  wire  _T_2 = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_2 ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_4 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_req_size; // @[Reg.scala 15:16]
  reg [86:0] r_req_user; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_9 = s3_io_isFinish ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_7 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_10 = s2_io_out_valid & s3_io_in_ready | _GEN_9; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_1_req_size; // @[Reg.scala 15:16]
  reg [86:0] r_1_req_user; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_0_tag; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_1_tag; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_2_tag; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_3_tag; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_3_data; // @[Reg.scala 15:16]
  reg  r_1_hit; // @[Reg.scala 15:16]
  reg [3:0] r_1_waymask; // @[Reg.scala 15:16]
  reg  r_1_mmio; // @[Reg.scala 15:16]
  reg  r_1_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] r_1_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] r_1_forwardData_waymask; // @[Reg.scala 15:16]
  CacheStage1 s1 ( // @[Cache.scala 484:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_user(s1_io_in_bits_user),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_user(s1_io_out_bits_req_user),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2 s2 ( // @[Cache.scala 485:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_user(s2_io_in_bits_req_user),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_user(s2_io_out_bits_req_user),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3 s3 ( // @[Cache.scala 486:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_user(s3_io_in_bits_req_user),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_out_bits_user(s3_io_out_bits_user),
    .io_isFinish(s3_io_isFinish),
    .io_flush(s3_io_flush),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 487:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 488:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_4 arb ( // @[Cache.scala 497:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_user(arb_io_in_0_bits_user),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_user(arb_io_out_bits_user)
  );
  assign io_in_req_ready = arb_io_in_0_ready; // @[Cache.scala 498:28]
  assign io_in_resp_valid = s3_io_out_valid; // @[Cache.scala 514:100]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 508:14]
  assign io_in_resp_bits_user = s3_io_out_bits_user; // @[Cache.scala 508:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 510:14]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 511:11]
  assign io_empty = ~s2_io_in_valid & ~s3_io_in_valid; // @[Cache.scala 512:31]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 500:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 500:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 500:12]
  assign s1_io_in_bits_user = arb_io_out_bits_user; // @[Cache.scala 500:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 532:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 533:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = r_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = r_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_user = r_req_user; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 539:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 542:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 541:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = r_1_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = r_1_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_user = r_1_req_user; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = r_1_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = r_1_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = r_1_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = r_1_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = r_1_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = r_1_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = r_1_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = r_1_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = r_1_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = r_1_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = r_1_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = r_1_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = r_1_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = r_1_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 508:14]
  assign s3_io_flush = io_flush[1]; // @[Cache.scala 509:26]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 534:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 510:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 511:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 511:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 511:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset | MOUFlushICache; // @[Cache.scala 494:37]
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 532:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 532:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 536:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 533:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 533:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 534:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 534:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 537:18]
  assign arb_io_in_0_valid = io_in_req_valid; // @[Cache.scala 498:28]
  assign arb_io_in_0_bits_addr = io_in_req_bits_addr; // @[Cache.scala 498:28]
  assign arb_io_in_0_bits_size = io_in_req_bits_size; // @[Cache.scala 498:28]
  assign arb_io_in_0_bits_user = io_in_req_bits_user; // @[Cache.scala 498:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 500:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_4) begin // @[Reg.scala 16:19]
      r_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_4) begin // @[Reg.scala 16:19]
      r_req_size <= s1_io_out_bits_req_size; // @[Reg.scala 16:23]
    end
    if (_T_4) begin // @[Reg.scala 16:19]
      r_req_user <= s1_io_out_bits_req_user; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[Pipeline.scala 27:20]
      REG_1 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_1 <= _GEN_10;
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_req_size <= s2_io_out_bits_req_size; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_req_user <= s2_io_out_bits_req_user; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_hit <= s2_io_out_bits_hit; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_req_size = _RAND_2[2:0];
  _RAND_3 = {3{`RANDOM}};
  r_req_user = _RAND_3[86:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_req_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_req_size = _RAND_6[2:0];
  _RAND_7 = {3{`RANDOM}};
  r_1_req_user = _RAND_7[86:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_metas_0_tag = _RAND_8[18:0];
  _RAND_9 = {1{`RANDOM}};
  r_1_metas_1_tag = _RAND_9[18:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_metas_2_tag = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  r_1_metas_3_tag = _RAND_11[18:0];
  _RAND_12 = {2{`RANDOM}};
  r_1_datas_0_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  r_1_datas_1_data = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  r_1_datas_2_data = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  r_1_datas_3_data = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_hit = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_waymask = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  r_1_mmio = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_1_isForwardData = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  r_1_forwardData_data_data = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  r_1_forwardData_waymask = _RAND_21[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SIMD_TLBEXEC_1(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_req_addr,
  input  [2:0]   io_in_bits_req_size,
  input  [3:0]   io_in_bits_req_cmd,
  input  [7:0]   io_in_bits_req_wmask,
  input  [63:0]  io_in_bits_req_wdata,
  input  [3:0]   io_in_bits_hitVec,
  input          io_in_bits_miss,
  input          io_in_bits_hitWB,
  input          io_in_bits_loadPF,
  input          io_in_bits_storePF,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_cmd,
  output [7:0]   io_out_bits_wmask,
  output [63:0]  io_out_bits_wdata,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_windex,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input          io_flush,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  input          io_pf_status_sum,
  input          io_pf_status_mxr,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output [38:0]  io_pf_addr,
  output         io_ipf,
  output         io_isFinish,
  input          ISAMO
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg  missLPF; // @[EmbeddedTLB.scala 687:24]
  reg  missSPF; // @[EmbeddedTLB.scala 688:24]
  wire [8:0] vpn_vpn0 = io_in_bits_req_addr[20:12]; // @[EmbeddedTLB.scala 694:54]
  wire [8:0] vpn_vpn1 = io_in_bits_req_addr[29:21]; // @[EmbeddedTLB.scala 694:54]
  wire [8:0] vpn_vpn2 = io_in_bits_req_addr[38:30]; // @[EmbeddedTLB.scala 694:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 696:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 696:30]
  wire  hit = io_in_valid & |io_in_bits_hitVec; // @[EmbeddedTLB.scala 701:25]
  wire  miss = io_in_valid & io_in_bits_miss; // @[EmbeddedTLB.scala 702:26]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_16 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_19 = {_T_16,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[EmbeddedTLB.scala 704:42]
  wire [3:0] waymask = hit ? io_in_bits_hitVec : victimWaymask; // @[EmbeddedTLB.scala 705:20]
  wire  _T_22 = io_in_bits_loadPF & io_in_valid; // @[EmbeddedTLB.scala 707:43]
  wire  _T_23 = io_in_bits_storePF & io_in_valid; // @[EmbeddedTLB.scala 708:45]
  wire  hitWB = io_in_bits_hitWB & io_in_valid; // @[EmbeddedTLB.scala 710:32]
  reg [2:0] state; // @[EmbeddedTLB.scala 733:22]
  wire  _T_107 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  reg  needFlush; // @[EmbeddedTLB.scala 746:26]
  wire  isFlush = needFlush | io_flush; // @[EmbeddedTLB.scala 748:27]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 741:49]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 741:49]
  wire [7:0] _T_98 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,
    memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 777:44]
  reg [1:0] level; // @[EmbeddedTLB.scala 734:22]
  wire  _T_110 = level == 2'h3; // @[EmbeddedTLB.scala 785:58]
  wire  _T_111 = level == 2'h2; // @[EmbeddedTLB.scala 785:73]
  wire  _T_122 = ~io_in_bits_req_cmd[0] & ~io_in_bits_req_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_124 = _T_122 & ~ISAMO; // @[EmbeddedTLB.scala 790:38]
  wire  _GEN_20 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? _T_122 & ~ISAMO : _T_22; // @[EmbeddedTLB.scala 786:60 790:22]
  wire  _T_165 = _T_98[0] & ~(io_pf_priviledgeMode == 2'h0 & ~_T_98[4]) & ~(io_pf_priviledgeMode == 2'h1 & _T_98[4] & ~
    io_pf_status_sum); // @[EmbeddedTLB.scala 804:87]
  wire  _T_169 = _T_165 & (_T_98[1] | io_pf_status_mxr & _T_98[3]); // @[EmbeddedTLB.scala 806:36]
  wire  _T_170 = _T_165 & _T_98[2]; // @[EmbeddedTLB.scala 807:37]
  wire  _T_175 = ~_T_98[6] | ~_T_98[7] & io_in_bits_req_cmd[0]; // @[EmbeddedTLB.scala 808:38]
  wire  _GEN_26 = ~_T_169 & _T_122 | ~_T_170 & io_in_bits_req_cmd[0] | _T_175 ? _T_124 : _T_22; // @[EmbeddedTLB.scala 821:92 823:22]
  wire  _GEN_34 = level != 2'h0 ? _GEN_26 : _T_22; // @[EmbeddedTLB.scala 803:36]
  wire  _GEN_42 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : _GEN_34; // @[EmbeddedTLB.scala 785:82]
  wire  _GEN_57 = isFlush ? _T_22 : _GEN_42; // @[EmbeddedTLB.scala 779:24]
  wire  _GEN_70 = _T_107 ? _GEN_57 : _T_22; // @[EmbeddedTLB.scala 778:33]
  wire  _GEN_124 = 3'h2 == state ? _GEN_70 : _T_22; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_138 = 3'h1 == state ? _T_22 : _GEN_124; // @[EmbeddedTLB.scala 753:18]
  wire  loadPF = 3'h0 == state ? _T_22 : _GEN_138; // @[EmbeddedTLB.scala 753:18]
  wire  _T_126 = io_in_bits_req_cmd[0] | ISAMO; // @[EmbeddedTLB.scala 792:40]
  wire  _GEN_22 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? io_in_bits_req_cmd[0] | ISAMO : _T_23; // @[EmbeddedTLB.scala 786:60 792:23]
  wire  _GEN_28 = ~_T_169 & _T_122 | ~_T_170 & io_in_bits_req_cmd[0] | _T_175 ? _T_126 : _T_23; // @[EmbeddedTLB.scala 821:92 825:23]
  wire  _GEN_36 = level != 2'h0 ? _GEN_28 : _T_23; // @[EmbeddedTLB.scala 803:36]
  wire  _GEN_44 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_22 : _GEN_36; // @[EmbeddedTLB.scala 785:82]
  wire  _GEN_58 = isFlush ? _T_23 : _GEN_44; // @[EmbeddedTLB.scala 779:24]
  wire  _GEN_71 = _T_107 ? _GEN_58 : _T_23; // @[EmbeddedTLB.scala 778:33]
  wire  _GEN_125 = 3'h2 == state ? _GEN_71 : _T_23; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_139 = 3'h1 == state ? _T_23 : _GEN_125; // @[EmbeddedTLB.scala 753:18]
  wire  storePF = 3'h0 == state ? _T_23 : _GEN_139; // @[EmbeddedTLB.scala 753:18]
  wire [120:0] _T_32 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_33 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_34 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_35 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_36 = _T_32 | _T_33; // @[Mux.scala 27:72]
  wire [120:0] _T_37 = _T_36 | _T_34; // @[Mux.scala 27:72]
  wire [120:0] _T_38 = _T_37 | _T_35; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_38[59:52]; // @[EmbeddedTLB.scala 718:70]
  wire [17:0] hitMeta_mask = _T_38[77:60]; // @[EmbeddedTLB.scala 718:70]
  wire [15:0] hitMeta_asid = _T_38[93:78]; // @[EmbeddedTLB.scala 718:70]
  wire [31:0] hitData_pteaddr = _T_38[31:0]; // @[EmbeddedTLB.scala 719:70]
  wire [19:0] hitData_ppn = _T_38[51:32]; // @[EmbeddedTLB.scala 719:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 720:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 720:38]
  wire [7:0] _T_69 = {io_in_bits_req_cmd[0],1'h1,6'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_70 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 723:79]
  wire [7:0] hitRefillFlag = _T_69 | _T_70; // @[EmbeddedTLB.scala 723:69]
  wire [39:0] _T_71 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 30:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 736:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 738:26]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 741:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 742:18]
  wire  _T_83 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[EmbeddedTLB.scala 746:26 749:{40,52}]
  wire  _GEN_4 = _T_83 & needFlush ? 1'h0 : _GEN_3; // @[EmbeddedTLB.scala 750:{37,49}]
  wire  _T_89 = ~isFlush; // @[EmbeddedTLB.scala 755:13]
  wire [31:0] _T_94 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 30:58]
  wire  _T_96 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_13 = _T_96 ? 3'h2 : state; // @[EmbeddedTLB.scala 733:22 773:{38,46}]
  wire  _GEN_15 = io_flush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 767:22 769:19]
  wire  _GEN_17 = io_flush ? 1'h0 : missSPF; // @[EmbeddedTLB.scala 767:22 771:17 688:24]
  wire  _GEN_18 = io_flush ? 1'h0 : missLPF; // @[EmbeddedTLB.scala 767:22 772:17 687:24]
  wire [8:0] _T_150 = _T_110 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 801:50]
  wire [31:0] _T_152 = {memRdata_ppn,_T_150,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_19 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? 3'h5 : 3'h1; // @[EmbeddedTLB.scala 786:60 787:73 800:19]
  wire  _GEN_21 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? loadPF : missLPF; // @[EmbeddedTLB.scala 786:60 791:23 687:24]
  wire  _GEN_23 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? storePF : missSPF; // @[EmbeddedTLB.scala 786:60 793:23 688:24]
  wire [31:0] _GEN_24 = ~_T_98[0] | ~_T_98[1] & _T_98[2] ? raddr : _T_152; // @[EmbeddedTLB.scala 742:18 786:60 801:19]
  wire [63:0] _T_177 = {56'h0,io_in_bits_req_cmd[0],7'h40}; // @[Cat.scala 30:58]
  wire [7:0] _T_180 = {_T_98[7],_T_98[6],_T_98[5],_T_98[4],_T_98[3],_T_98[2],_T_98[1],_T_98[0]}; // @[EmbeddedTLB.scala 810:79]
  wire [7:0] _T_181 = _T_69 | _T_180; // @[EmbeddedTLB.scala 810:68]
  wire [63:0] _T_182 = io_mem_resp_bits_rdata | _T_177; // @[EmbeddedTLB.scala 811:50]
  wire [2:0] _GEN_25 = ~_T_169 & _T_122 | ~_T_170 & io_in_bits_req_cmd[0] | _T_175 ? 3'h5 : 3'h4; // @[EmbeddedTLB.scala 821:92 822:21 828:21]
  wire  _GEN_27 = ~_T_169 & _T_122 | ~_T_170 & io_in_bits_req_cmd[0] | _T_175 ? loadPF : missLPF; // @[EmbeddedTLB.scala 821:92 824:23 687:24]
  wire  _GEN_29 = ~_T_169 & _T_122 | ~_T_170 & io_in_bits_req_cmd[0] | _T_175 ? storePF : missSPF; // @[EmbeddedTLB.scala 821:92 826:23 688:24]
  wire  _GEN_30 = ~_T_169 & _T_122 | ~_T_170 & io_in_bits_req_cmd[0] | _T_175 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 821:92 829:30]
  wire [17:0] _T_206 = _T_111 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 832:59]
  wire [17:0] _T_207 = _T_110 ? 18'h0 : _T_206; // @[EmbeddedTLB.scala 832:26]
  wire [7:0] _GEN_31 = level != 2'h0 ? _T_181 : 8'h0; // @[EmbeddedTLB.scala 803:36 810:26]
  wire [63:0] _GEN_32 = level != 2'h0 ? _T_182 : memRespStore; // @[EmbeddedTLB.scala 803:36 811:24 736:25]
  wire [2:0] _GEN_33 = level != 2'h0 ? _GEN_25 : state; // @[EmbeddedTLB.scala 733:22 803:36]
  wire  _GEN_35 = level != 2'h0 ? _GEN_27 : missLPF; // @[EmbeddedTLB.scala 687:24 803:36]
  wire  _GEN_37 = level != 2'h0 ? _GEN_29 : missSPF; // @[EmbeddedTLB.scala 688:24 803:36]
  wire  _GEN_38 = level != 2'h0 & _GEN_30; // @[EmbeddedTLB.scala 803:36]
  wire [17:0] _GEN_39 = level != 2'h0 ? _T_207 : 18'h3ffff; // @[EmbeddedTLB.scala 803:36 832:20]
  wire [17:0] _GEN_50 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_39; // @[EmbeddedTLB.scala 785:82]
  wire [17:0] _GEN_63 = isFlush ? 18'h3ffff : _GEN_50; // @[EmbeddedTLB.scala 779:24]
  wire [17:0] _GEN_76 = _T_107 ? _GEN_63 : 18'h3ffff; // @[EmbeddedTLB.scala 778:33]
  wire [17:0] _GEN_130 = 3'h2 == state ? _GEN_76 : 18'h3ffff; // @[EmbeddedTLB.scala 753:18]
  wire [17:0] _GEN_144 = 3'h1 == state ? 18'h3ffff : _GEN_130; // @[EmbeddedTLB.scala 753:18]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_144; // @[EmbeddedTLB.scala 753:18]
  wire [17:0] _GEN_40 = level != 2'h0 ? missMask : missMaskStore; // @[EmbeddedTLB.scala 803:36 833:25 738:26]
  wire [2:0] _GEN_41 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_33; // @[EmbeddedTLB.scala 785:82]
  wire  _GEN_43 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_21 : _GEN_35; // @[EmbeddedTLB.scala 785:82]
  wire  _GEN_45 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_23 : _GEN_37; // @[EmbeddedTLB.scala 785:82]
  wire [31:0] _GEN_46 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_24 : raddr; // @[EmbeddedTLB.scala 742:18 785:82]
  wire [7:0] _GEN_47 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_31; // @[EmbeddedTLB.scala 785:82]
  wire [63:0] _GEN_48 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_32; // @[EmbeddedTLB.scala 736:25 785:82]
  wire  _GEN_49 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_38; // @[EmbeddedTLB.scala 785:82]
  wire [17:0] _GEN_51 = ~(_T_98[1] | _T_98[3]) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_40; // @[EmbeddedTLB.scala 738:26 785:82]
  wire [2:0] _GEN_52 = isFlush ? 3'h0 : _GEN_41; // @[EmbeddedTLB.scala 779:24 780:17]
  wire  _GEN_54 = isFlush ? 1'h0 : _GEN_45; // @[EmbeddedTLB.scala 779:24 782:19]
  wire  _GEN_55 = isFlush ? 1'h0 : _GEN_43; // @[EmbeddedTLB.scala 779:24 783:19]
  wire  _GEN_56 = isFlush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 779:24 784:21]
  wire [31:0] _GEN_59 = isFlush ? raddr : _GEN_46; // @[EmbeddedTLB.scala 742:18 779:24]
  wire [7:0] _GEN_60 = isFlush ? 8'h0 : _GEN_47; // @[EmbeddedTLB.scala 779:24]
  wire [63:0] _GEN_61 = isFlush ? memRespStore : _GEN_48; // @[EmbeddedTLB.scala 779:24 736:25]
  wire  _GEN_62 = isFlush ? 1'h0 : _GEN_49; // @[EmbeddedTLB.scala 779:24]
  wire [17:0] _GEN_64 = isFlush ? missMaskStore : _GEN_51; // @[EmbeddedTLB.scala 779:24 738:26]
  wire [1:0] _T_209 = level - 2'h1; // @[EmbeddedTLB.scala 835:24]
  wire [2:0] _GEN_65 = _T_107 ? _GEN_52 : state; // @[EmbeddedTLB.scala 733:22 778:33]
  wire  _GEN_67 = _T_107 ? _GEN_54 : missSPF; // @[EmbeddedTLB.scala 688:24 778:33]
  wire  _GEN_68 = _T_107 ? _GEN_55 : missLPF; // @[EmbeddedTLB.scala 687:24 778:33]
  wire  _GEN_69 = _T_107 ? _GEN_56 : _GEN_4; // @[EmbeddedTLB.scala 778:33]
  wire [7:0] _GEN_73 = _T_107 ? _GEN_60 : 8'h0; // @[EmbeddedTLB.scala 778:33]
  wire  _GEN_75 = _T_107 & _GEN_62; // @[EmbeddedTLB.scala 778:33]
  wire [1:0] _GEN_78 = _T_107 ? _T_209 : level; // @[EmbeddedTLB.scala 778:33 835:15 734:22]
  wire [2:0] _GEN_79 = _T_96 ? 3'h6 : state; // @[EmbeddedTLB.scala 733:22 846:{38,46}]
  wire [2:0] _GEN_80 = io_flush ? 3'h0 : _GEN_79; // @[EmbeddedTLB.scala 840:22 841:15]
  wire [2:0] _GEN_81 = isFlush ? 3'h0 : 3'h4; // @[EmbeddedTLB.scala 851:22 852:17 858:17]
  wire  _GEN_82 = isFlush ? 1'h0 : missSPF; // @[EmbeddedTLB.scala 851:22 855:19 688:24]
  wire  _GEN_83 = isFlush ? 1'h0 : missLPF; // @[EmbeddedTLB.scala 851:22 856:19 687:24]
  wire [2:0] _GEN_84 = _T_107 ? _GEN_81 : state; // @[EmbeddedTLB.scala 733:22 850:32]
  wire  _GEN_87 = _T_107 ? _GEN_82 : missSPF; // @[EmbeddedTLB.scala 688:24 850:32]
  wire  _GEN_88 = _T_107 ? _GEN_83 : missLPF; // @[EmbeddedTLB.scala 687:24 850:32]
  wire [2:0] _GEN_89 = _T_83 | io_flush ? 3'h0 : state; // @[EmbeddedTLB.scala 863:56 864:13 733:22]
  wire  _GEN_91 = _T_83 | io_flush ? 1'h0 : missSPF; // @[EmbeddedTLB.scala 863:56 866:15 688:24]
  wire  _GEN_92 = _T_83 | io_flush ? 1'h0 : missLPF; // @[EmbeddedTLB.scala 863:56 867:15 687:24]
  wire  _GEN_93 = _T_83 | io_flush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 863:56 868:17]
  wire [2:0] _GEN_99 = 3'h5 == state ? _GEN_89 : state; // @[EmbeddedTLB.scala 753:18 733:22]
  wire  _GEN_100 = 3'h5 == state ? _GEN_91 : missSPF; // @[EmbeddedTLB.scala 753:18 688:24]
  wire  _GEN_101 = 3'h5 == state ? _GEN_92 : missLPF; // @[EmbeddedTLB.scala 753:18 687:24]
  wire  _GEN_103 = 3'h5 == state ? _GEN_93 : _GEN_4; // @[EmbeddedTLB.scala 753:18]
  wire [2:0] _GEN_104 = 3'h4 == state ? _GEN_89 : _GEN_99; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_106 = 3'h4 == state ? _GEN_91 : _GEN_100; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_107 = 3'h4 == state ? _GEN_92 : _GEN_101; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_108 = 3'h4 == state ? _GEN_93 : _GEN_103; // @[EmbeddedTLB.scala 753:18]
  wire [2:0] _GEN_109 = 3'h6 == state ? _GEN_84 : _GEN_104; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_110 = 3'h6 == state ? _GEN_69 : _GEN_108; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_112 = 3'h6 == state ? _GEN_87 : _GEN_106; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_113 = 3'h6 == state ? _GEN_88 : _GEN_107; // @[EmbeddedTLB.scala 753:18]
  wire [2:0] _GEN_114 = 3'h3 == state ? _GEN_80 : _GEN_109; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_115 = 3'h3 == state ? _GEN_15 : _GEN_110; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_117 = 3'h3 == state ? _GEN_17 : _GEN_112; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_118 = 3'h3 == state ? _GEN_18 : _GEN_113; // @[EmbeddedTLB.scala 753:18]
  wire [7:0] _GEN_127 = 3'h2 == state ? _GEN_73 : 8'h0; // @[EmbeddedTLB.scala 753:18]
  wire [7:0] _GEN_141 = 3'h1 == state ? 8'h0 : _GEN_127; // @[EmbeddedTLB.scala 753:18]
  wire  _GEN_143 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_75; // @[EmbeddedTLB.scala 753:18]
  wire [7:0] missRefillFlag = 3'h0 == state ? 8'h0 : _GEN_141; // @[EmbeddedTLB.scala 753:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_143; // @[EmbeddedTLB.scala 753:18]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 883:23]
  wire [31:0] _T_221 = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 884:35]
  wire  _T_226 = ~io_flush; // @[EmbeddedTLB.scala 885:77]
  wire [15:0] _T_240 = hitWB ? hitMeta_asid : satp_asid; // @[EmbeddedTLB.scala 891:15]
  wire [17:0] _T_241 = hitWB ? hitMeta_mask : missMask; // @[EmbeddedTLB.scala 891:59]
  wire [7:0] _T_242 = hitWB ? hitRefillFlag : missRefillFlag; // @[EmbeddedTLB.scala 892:15]
  wire [19:0] _T_243 = hitWB ? hitData_ppn : memRdata_ppn; // @[EmbeddedTLB.scala 892:64]
  wire [59:0] lo_5 = {_T_242,_T_243,_T_221}; // @[Cat.scala 30:58]
  wire [60:0] hi_8 = {vpn_vpn2,vpn_vpn1,vpn_vpn0,_T_240,_T_241}; // @[Cat.scala 30:58]
  wire [31:0] _T_247 = {hitData_ppn,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_249 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_250 = _T_247 & _T_249; // @[BitUtils.scala 32:13]
  wire [31:0] _T_251 = ~_T_249; // @[BitUtils.scala 32:38]
  wire [31:0] _T_252 = io_in_bits_req_addr[31:0] & _T_251; // @[BitUtils.scala 32:36]
  wire [31:0] _T_253 = _T_250 | _T_252; // @[BitUtils.scala 32:25]
  wire [31:0] _T_266 = {memRespStore[29:10],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_268 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_269 = _T_266 & _T_268; // @[BitUtils.scala 32:13]
  wire [31:0] _T_270 = ~_T_268; // @[BitUtils.scala 32:38]
  wire [31:0] _T_271 = io_in_bits_req_addr[31:0] & _T_270; // @[BitUtils.scala 32:36]
  wire [31:0] _T_272 = _T_269 | _T_271; // @[BitUtils.scala 32:25]
  wire  _T_276 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 176:23]
  assign io_in_ready = ~io_in_valid | _T_83 & io_mdReady; // @[EmbeddedTLB.scala 900:31]
  assign io_out_valid = _T_226 & io_in_valid & (state == 3'h4 & ~(_T_276 | loadPF | storePF | missLPF | missSPF | io_ipf
    )); // @[EmbeddedTLB.scala 898:43]
  assign io_out_bits_addr = hit ? _T_253 : _T_272; // @[EmbeddedTLB.scala 897:26]
  assign io_out_bits_size = io_in_bits_req_size; // @[EmbeddedTLB.scala 896:15]
  assign io_out_bits_cmd = io_in_bits_req_cmd; // @[EmbeddedTLB.scala 896:15]
  assign io_out_bits_wmask = io_in_bits_req_wmask; // @[EmbeddedTLB.scala 896:15]
  assign io_out_bits_wdata = io_in_bits_req_wdata; // @[EmbeddedTLB.scala 896:15]
  assign io_mdWrite_wen = io_in_valid & (missMetaRefill & _T_89 | hitWB & state == 3'h0 & _T_89); // @[EmbeddedTLB.scala 889:38]
  assign io_mdWrite_windex = io_in_bits_req_addr[15:12]; // @[TLB.scala 200:19]
  assign io_mdWrite_waymask = hit ? io_in_bits_hitVec : victimWaymask; // @[EmbeddedTLB.scala 705:20]
  assign io_mdWrite_wdata = {hi_8,lo_5}; // @[Cat.scala 30:58]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~io_flush; // @[EmbeddedTLB.scala 885:74]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 884:35]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[EmbeddedTLB.scala 884:138]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 886:21]
  assign io_pf_loadPF = (loadPF | missLPF) & io_in_valid; // @[EmbeddedTLB.scala 713:39]
  assign io_pf_storePF = (storePF | missSPF) & io_in_valid; // @[EmbeddedTLB.scala 714:41]
  assign io_pf_addr = io_in_bits_req_addr; // @[EmbeddedTLB.scala 715:14]
  assign io_ipf = 1'h0; // @[EmbeddedTLB.scala 902:16]
  assign io_isFinish = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  always @(posedge clock) begin
    if (reset) begin // @[EmbeddedTLB.scala 687:24]
      missLPF <= 1'h0; // @[EmbeddedTLB.scala 687:24]
    end else if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
        if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
          missLPF <= 1'h0; // @[EmbeddedTLB.scala 772:17]
        end
      end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        missLPF <= _GEN_68;
      end else begin
        missLPF <= _GEN_118;
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 688:24]
      missSPF <= 1'h0; // @[EmbeddedTLB.scala 688:24]
    end else if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
        if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
          missSPF <= 1'h0; // @[EmbeddedTLB.scala 771:17]
        end
      end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        missSPF <= _GEN_67;
      end else begin
        missSPF <= _GEN_117;
      end
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_19;
    end
    if (reset) begin // @[EmbeddedTLB.scala 733:22]
      state <= 3'h0; // @[EmbeddedTLB.scala 733:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (~isFlush & hitWB) begin // @[EmbeddedTLB.scala 755:32]
        state <= 3'h3; // @[EmbeddedTLB.scala 756:15]
      end else if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
        state <= 3'h1; // @[EmbeddedTLB.scala 759:15]
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
        state <= 3'h0; // @[EmbeddedTLB.scala 768:15]
      end else begin
        state <= _GEN_13;
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
      state <= _GEN_65;
    end else begin
      state <= _GEN_114;
    end
    if (reset) begin // @[EmbeddedTLB.scala 746:26]
      needFlush <= 1'h0; // @[EmbeddedTLB.scala 746:26]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (~isFlush & hitWB) begin // @[EmbeddedTLB.scala 755:32]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 757:19]
      end else if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 762:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (io_flush) begin // @[EmbeddedTLB.scala 767:22]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 769:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
      needFlush <= _GEN_69;
    end else begin
      needFlush <= _GEN_115;
    end
    if (reset) begin // @[EmbeddedTLB.scala 734:22]
      level <= 2'h3; // @[EmbeddedTLB.scala 734:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (!(~isFlush & hitWB)) begin // @[EmbeddedTLB.scala 755:32]
        if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
          level <= 2'h3; // @[EmbeddedTLB.scala 761:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        level <= _GEN_78;
      end
    end
    if (hitWB) begin // @[Reg.scala 16:19]
      hitWBStore <= _T_71; // @[Reg.scala 16:23]
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
          if (_T_107) begin // @[EmbeddedTLB.scala 778:33]
            memRespStore <= _GEN_61;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
          if (_T_107) begin // @[EmbeddedTLB.scala 778:33]
            missMaskStore <= _GEN_64;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[EmbeddedTLB.scala 753:18]
      if (!(~isFlush & hitWB)) begin // @[EmbeddedTLB.scala 755:32]
        if (miss & _T_89) begin // @[EmbeddedTLB.scala 758:37]
          raddr <= _T_94; // @[EmbeddedTLB.scala 760:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 753:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 753:18]
        if (_T_107) begin // @[EmbeddedTLB.scala 778:33]
          raddr <= _GEN_59;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  missLPF = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  missSPF = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  REG = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  needFlush = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  level = _RAND_5[1:0];
  _RAND_6 = {2{`RANDOM}};
  hitWBStore = _RAND_6[39:0];
  _RAND_7 = {2{`RANDOM}};
  memRespStore = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  missMaskStore = _RAND_8[17:0];
  _RAND_9 = {1{`RANDOM}};
  raddr = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBEmpty_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  wire  _T_1 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = ~io_in_valid | _T_1; // @[EmbeddedTLB.scala 407:31]
  assign io_out_valid = io_in_valid; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 406:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_windex,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  input  [3:0]   io_rindex,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_0_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_0_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_1 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_1_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_1_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_2 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_2_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_2_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_3 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_3_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_3_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg  resetState; // @[EmbeddedTLB.scala 55:27]
  reg [3:0] resetSet; // @[Counter.scala 60:40]
  wire  wrap_wrap = resetSet == 4'hf; // @[Counter.scala 72:24]
  wire [3:0] _wrap_value_T_1 = resetSet + 4'h1; // @[Counter.scala 76:24]
  wire  resetFinish = resetState & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[EmbeddedTLB.scala 57:22 55:27 57:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 66:20]
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = io_rindex;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = io_rindex;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = io_rindex;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = io_rindex;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 72:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    resetState <= reset | _GEN_2; // @[EmbeddedTLB.scala 55:{27,27}]
    if (reset) begin // @[Counter.scala 60:40]
      resetSet <= 4'h0; // @[Counter.scala 60:40]
    end else if (resetState) begin // @[Counter.scala 118:17]
      resetSet <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SIMD_TLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_flush,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_csrMMU_status_sum,
  input         io_csrMMU_status_mxr,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  output [38:0] io_csrMMU_addr,
  output        _T_408_0,
  input  [63:0] CSRSATP,
  output        ismmio_0,
  input         ISAMO,
  output        vmEnable_0,
  output        _T_407_0,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 443:23]
  wire [38:0] tlbExec_io_in_bits_req_addr; // @[EmbeddedTLB.scala 443:23]
  wire [2:0] tlbExec_io_in_bits_req_size; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_in_bits_req_cmd; // @[EmbeddedTLB.scala 443:23]
  wire [7:0] tlbExec_io_in_bits_req_wmask; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_in_bits_req_wdata; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_in_bits_hitVec; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_miss; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_hitWB; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_loadPF; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_in_bits_storePF; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 443:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 443:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[EmbeddedTLB.scala 443:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 443:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 443:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 443:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_flush; // @[EmbeddedTLB.scala 443:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 443:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_pf_status_sum; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_pf_status_mxr; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 443:23]
  wire [38:0] tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 443:23]
  wire  tlbExec_ISAMO; // @[EmbeddedTLB.scala 443:23]
  wire  tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 444:24]
  wire  tlbEmpty_io_in_valid; // @[EmbeddedTLB.scala 444:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[EmbeddedTLB.scala 444:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[EmbeddedTLB.scala 444:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[EmbeddedTLB.scala 444:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[EmbeddedTLB.scala 444:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[EmbeddedTLB.scala 444:24]
  wire  tlbEmpty_io_out_ready; // @[EmbeddedTLB.scala 444:24]
  wire  tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 444:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 444:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 444:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 444:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 444:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 444:24]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 445:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 445:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 445:21]
  wire [3:0] mdTLB_io_write_windex; // @[EmbeddedTLB.scala 445:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 445:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 445:21]
  wire [3:0] mdTLB_io_rindex; // @[EmbeddedTLB.scala 445:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 445:21]
  reg  REG; // @[EmbeddedTLB.scala 454:30]
  reg  REG_1; // @[EmbeddedTLB.scala 455:31]
  reg [38:0] REG_2; // @[EmbeddedTLB.scala 456:28]
  reg [120:0] r__0; // @[Reg.scala 15:16]
  reg [120:0] r__1; // @[Reg.scala 15:16]
  reg [120:0] r__2; // @[Reg.scala 15:16]
  reg [120:0] r__3; // @[Reg.scala 15:16]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 470:57]
  wire [120:0] _WIRE_46 = mdTLB_io_tlbmd_3;
  wire [26:0] _T_208 = {9'h1ff,_WIRE_46[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_209 = _T_208 & _WIRE_46[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_207 = {io_in_req_bits_addr[38:30],io_in_req_bits_addr[29:21],io_in_req_bits_addr[20:12]}; // @[EmbeddedTLB.scala 531:224]
  wire [26:0] _T_211 = _T_208 & _T_207; // @[TLB.scala 131:84]
  wire  _T_212 = _T_209 == _T_211; // @[TLB.scala 131:48]
  wire  _T_213 = _WIRE_46[52] & _WIRE_46[93:78] == CSRSATP[59:44] & _T_212; // @[EmbeddedTLB.scala 531:155]
  wire [120:0] _WIRE_34 = mdTLB_io_tlbmd_2;
  wire [26:0] _T_163 = {9'h1ff,_WIRE_34[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_164 = _T_163 & _WIRE_34[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_166 = _T_163 & _T_207; // @[TLB.scala 131:84]
  wire  _T_167 = _T_164 == _T_166; // @[TLB.scala 131:48]
  wire  _T_168 = _WIRE_34[52] & _WIRE_34[93:78] == CSRSATP[59:44] & _T_167; // @[EmbeddedTLB.scala 531:155]
  wire [120:0] _WIRE_22 = mdTLB_io_tlbmd_1;
  wire [26:0] _T_118 = {9'h1ff,_WIRE_22[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_119 = _T_118 & _WIRE_22[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_121 = _T_118 & _T_207; // @[TLB.scala 131:84]
  wire  _T_122 = _T_119 == _T_121; // @[TLB.scala 131:48]
  wire  _T_123 = _WIRE_22[52] & _WIRE_22[93:78] == CSRSATP[59:44] & _T_122; // @[EmbeddedTLB.scala 531:155]
  wire [120:0] _WIRE_10 = mdTLB_io_tlbmd_0;
  wire [26:0] _T_73 = {9'h1ff,_WIRE_10[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_74 = _T_73 & _WIRE_10[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_76 = _T_73 & _T_207; // @[TLB.scala 131:84]
  wire  _T_77 = _T_74 == _T_76; // @[TLB.scala 131:48]
  wire  _T_78 = _WIRE_10[52] & _WIRE_10[93:78] == CSRSATP[59:44] & _T_77; // @[EmbeddedTLB.scala 531:155]
  wire [3:0] _T_214 = {_T_213,_T_168,_T_123,_T_78}; // @[EmbeddedTLB.scala 531:234]
  wire  _T_217 = |_T_214; // @[EmbeddedTLB.scala 533:43]
  wire  _T_219 = io_in_req_valid & ~(|_T_214); // @[EmbeddedTLB.scala 533:32]
  wire  _T_216 = io_in_req_valid & _T_217; // @[EmbeddedTLB.scala 532:31]
  reg [63:0] REG_5; // @[LFSR64.scala 25:23]
  wire [3:0] _T_232 = 4'h1 << REG_5[1:0]; // @[EmbeddedTLB.scala 535:44]
  wire [3:0] _T_233 = _T_216 ? _T_214 : _T_232; // @[EmbeddedTLB.scala 536:22]
  wire [120:0] _T_238 = _T_233[0] ? mdTLB_io_tlbmd_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_239 = _T_233[1] ? mdTLB_io_tlbmd_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_242 = _T_238 | _T_239; // @[Mux.scala 27:72]
  wire [120:0] _T_240 = _T_233[2] ? mdTLB_io_tlbmd_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_243 = _T_242 | _T_240; // @[Mux.scala 27:72]
  wire [120:0] _T_241 = _T_233[3] ? mdTLB_io_tlbmd_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_244 = _T_243 | _T_241; // @[Mux.scala 27:72]
  wire  _T_303 = _T_216 & ~(io_csrMMU_priviledgeMode == 2'h0 & ~_T_244[56]) & ~(io_csrMMU_priviledgeMode == 2'h1 &
    _T_244[56] & ~io_csrMMU_status_sum); // @[EmbeddedTLB.scala 557:96]
  wire  _T_307 = _T_303 & (_T_244[53] | io_csrMMU_status_mxr & _T_244[55]); // @[EmbeddedTLB.scala 559:28]
  wire  _T_314 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_316 = ~_T_307 & _T_314 & _T_216; // @[EmbeddedTLB.scala 572:42]
  wire  _T_318 = ~_T_307 & _T_314 & _T_216 & ~ISAMO; // @[EmbeddedTLB.scala 572:49]
  wire  _T_308 = _T_303 & _T_244[54]; // @[EmbeddedTLB.scala 560:29]
  wire  _T_332 = ~_T_308 & io_in_req_bits_cmd[0] & _T_216 | _T_316 & ISAMO; // @[EmbeddedTLB.scala 573:54]
  wire  _T_283 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 176:23]
  wire  _T_286 = _T_216 & (~_T_244[58] | ~_T_244[59] & io_in_req_bits_cmd[0]) & ~(_T_318 | _T_332 | _T_283); // @[EmbeddedTLB.scala 552:83]
  wire  _T_374 = _T_219 | _T_286 | _T_318 | _T_332; // @[EmbeddedTLB.scala 609:75]
  wire  tlbexec_inbundle_valid = ~vmEnable ? 1'h0 : io_in_req_valid & (_T_219 | _T_286 | _T_318 | _T_332); // @[EmbeddedTLB.scala 507:19 508:28 609:28]
  wire  mdUpdate = tlbexec_inbundle_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 482:26]
  reg  REG_3; // @[EmbeddedTLB.scala 473:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : REG_3; // @[EmbeddedTLB.scala 473:24 474:{25,33}]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[EmbeddedTLB.scala 475:{50,58}]
  reg [38:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_1_req_size; // @[Reg.scala 15:16]
  reg [3:0] r_1_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_1_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_1_req_wdata; // @[Reg.scala 15:16]
  reg [3:0] r_1_hitVec; // @[Reg.scala 15:16]
  reg  r_1_miss; // @[Reg.scala 15:16]
  reg  r_1_hitWB; // @[Reg.scala 15:16]
  reg  r_1_loadPF; // @[Reg.scala 15:16]
  reg  r_1_storePF; // @[Reg.scala 15:16]
  wire  _T_15 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG_4; // @[Pipeline.scala 24:24]
  wire  _GEN_18 = _T_15 ? 1'h0 : REG_4; // @[Pipeline.scala 24:24 25:{25,33}]
  reg  state; // @[EmbeddedTLB.scala 505:22]
  wire  _T_333 = ~state; // @[EmbeddedTLB.scala 577:32]
  wire  _T_341 = ~state ? _T_216 & ~_T_286 & ~(_T_283 | _T_318 | _T_332) : tlbExec_io_out_valid; // @[EmbeddedTLB.scala 577:25]
  wire  out_req_valid = ~vmEnable ? 1'h0 : _T_341; // @[EmbeddedTLB.scala 507:19 521:19 577:19]
  wire  _T_16 = out_req_valid & tlbEmpty_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_19 = out_req_valid & tlbEmpty_io_in_ready | _GEN_18; // @[Pipeline.scala 26:{38,46}]
  reg [38:0] r_2_addr; // @[Reg.scala 15:16]
  reg [2:0] r_2_size; // @[Reg.scala 15:16]
  reg [3:0] r_2_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_2_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_2_wdata; // @[Reg.scala 15:16]
  wire [31:0] _T_344 = {_T_244[51:32],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_346 = {2'h3,_T_244[77:60],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_347 = _T_344 & _T_346; // @[BitUtils.scala 32:13]
  wire [31:0] _T_348 = ~_T_346; // @[BitUtils.scala 32:38]
  wire [31:0] _T_349 = io_in_req_bits_addr[31:0] & _T_348; // @[BitUtils.scala 32:36]
  wire [31:0] _T_350 = _T_347 | _T_349; // @[BitUtils.scala 32:25]
  wire [31:0] _T_351 = _T_333 ? _T_350 : tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 578:29]
  wire [31:0] _GEN_57 = ~vmEnable ? tlbExec_io_out_bits_addr : _T_351; // @[EmbeddedTLB.scala 495:16 507:19 578:23]
  wire [38:0] out_req_bits_addr = {{7'd0}, _GEN_57}; // @[EmbeddedTLB.scala 494:21]
  wire  _T_20 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_22 = io_out_req_bits_addr < 32'h40000000; // @[NutCore.scala 92:35]
  wire  _T_26 = io_out_req_bits_addr >= 32'h40600000 & io_out_req_bits_addr < 32'h41600000; // @[NutCore.scala 92:26]
  wire  _T_27 = _T_22 | _T_26; // @[NutCore.scala 93:15]
  wire  _T_226 = REG_5[0] ^ REG_5[1] ^ REG_5[3] ^ REG_5[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_229 = {_T_226,REG_5[63:1]}; // @[Cat.scala 30:58]
  wire  out_req_ready = ~vmEnable ? 1'h0 : tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 507:19 522:19 Pipeline.scala 29:16]
  wire  _T_352 = out_req_ready & out_req_valid; // @[Decoupled.scala 40:37]
  wire  tlbexec_inbundle_ready = tlbExec_io_in_ready; // @[EmbeddedTLB.scala 478:16 490:30]
  wire  _T_361 = tlbexec_inbundle_ready & tlbexec_inbundle_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_374 & ~io_flush & _T_361 | state; // @[EmbeddedTLB.scala 588:105 589:17 505:22]
  wire  _GEN_30 = _T_352 | io_flush ? 1'h0 : state; // @[EmbeddedTLB.scala 593:41 595:17 505:22]
  wire  _GEN_31 = ~io_in_req_valid ? 1'h0 : _GEN_30; // @[EmbeddedTLB.scala 597:31 598:17]
  wire  _GEN_32 = ~io_in_req_valid | io_flush; // @[EmbeddedTLB.scala 448:20 597:31 599:28]
  wire  _GEN_34 = state ? _GEN_32 : io_flush; // @[EmbeddedTLB.scala 586:19 448:20]
  wire  _GEN_36 = _T_333 ? io_flush : _GEN_34; // @[EmbeddedTLB.scala 586:19 448:20]
  wire  _T_394 = out_req_bits_addr < 39'h40000000; // @[NutCore.scala 92:35]
  wire  _T_398 = out_req_bits_addr >= 39'h40600000 & out_req_bits_addr < 39'h41600000; // @[NutCore.scala 92:26]
  wire  _T_399 = _T_394 | _T_398; // @[NutCore.scala 93:15]
  wire  _T_406 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[Bundle.scala 176:23]
  wire  _T_407 = _T_352 | _T_406; // @[EmbeddedTLB.scala 627:38]
  wire  _T_408 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 176:23]
  wire  ismmio = ~vmEnable ? _T_20 & _T_27 : _T_352 & _T_399; // @[EmbeddedTLB.scala 507:19 523:12 618:12]
  SIMD_TLBEXEC_1 tlbExec ( // @[EmbeddedTLB.scala 443:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_req_addr(tlbExec_io_in_bits_req_addr),
    .io_in_bits_req_size(tlbExec_io_in_bits_req_size),
    .io_in_bits_req_cmd(tlbExec_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(tlbExec_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(tlbExec_io_in_bits_req_wdata),
    .io_in_bits_hitVec(tlbExec_io_in_bits_hitVec),
    .io_in_bits_miss(tlbExec_io_in_bits_miss),
    .io_in_bits_hitWB(tlbExec_io_in_bits_hitWB),
    .io_in_bits_loadPF(tlbExec_io_in_bits_loadPF),
    .io_in_bits_storePF(tlbExec_io_in_bits_storePF),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_addr(tlbExec_io_pf_addr),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish),
    .ISAMO(tlbExec_ISAMO)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[EmbeddedTLB.scala 444:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[EmbeddedTLB.scala 445:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : _T_352; // @[EmbeddedTLB.scala 507:19 513:21 580:21]
  assign io_in_resp_valid = io_out_resp_valid; // @[EmbeddedTLB.scala 620:14]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 620:14]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 501:18 507:19 512:22]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 501:18 507:19 514:26]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 501:18 507:19 515:26]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 501:18 507:19 516:25]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 501:18 507:19 517:27]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 501:18 507:19 518:27]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 450:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 450:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 450:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 450:18]
  assign io_csrMMU_loadPF = REG; // @[EmbeddedTLB.scala 454:20]
  assign io_csrMMU_storePF = REG_1; // @[EmbeddedTLB.scala 455:21]
  assign io_csrMMU_addr = REG_2; // @[EmbeddedTLB.scala 456:18]
  assign _T_408_0 = _T_283;
  assign ismmio_0 = ismmio;
  assign vmEnable_0 = vmEnable;
  assign _T_407_0 = _T_407;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = REG_3; // @[EmbeddedTLB.scala 480:17]
  assign tlbExec_io_in_bits_req_addr = r_1_req_addr; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_req_size = r_1_req_size; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_req_cmd = r_1_req_cmd; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_req_wmask = r_1_req_wmask; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_req_wdata = r_1_req_wdata; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_hitVec = r_1_hitVec; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_miss = r_1_miss; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_hitWB = r_1_hitWB; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_loadPF = r_1_loadPF; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_in_bits_storePF = r_1_storePF; // @[EmbeddedTLB.scala 479:16]
  assign tlbExec_io_out_ready = ~vmEnable | _T_352; // @[EmbeddedTLB.scala 507:19 509:26 579:26]
  assign tlbExec_io_md_0 = r__0; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_md_1 = r__1; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_md_2 = r__2; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_md_3 = r__3; // @[EmbeddedTLB.scala 457:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 458:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 450:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 450:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 450:18]
  assign tlbExec_io_flush = ~vmEnable ? io_flush : _GEN_36; // @[EmbeddedTLB.scala 507:19 448:20]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 449:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 451:32]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[EmbeddedTLB.scala 452:28]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 453:28]
  assign tlbExec_ISAMO = ISAMO;
  assign tlbEmpty_io_in_valid = REG_4; // @[Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = r_2_addr[31:0]; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = r_2_size; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = r_2_cmd; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = r_2_wmask; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = r_2_wdata; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[EmbeddedTLB.scala 501:18 507:19 511:52]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 467:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 460:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 460:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 460:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 460:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[TLB.scala 200:19]
  always @(posedge clock) begin
    REG <= tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 454:30]
    REG_1 <= tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 455:31]
    REG_2 <= tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 456:28]
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__0 <= mdTLB_io_tlbmd_0; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__1 <= mdTLB_io_tlbmd_1; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__2 <= mdTLB_io_tlbmd_2; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__3 <= mdTLB_io_tlbmd_3; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG_5 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG_5 == 64'h0) begin // @[LFSR64.scala 28:18]
      REG_5 <= 64'h1;
    end else begin
      REG_5 <= _T_229;
    end
    if (reset) begin // @[EmbeddedTLB.scala 473:24]
      REG_3 <= 1'h0; // @[EmbeddedTLB.scala 473:24]
    end else if (io_flush) begin // @[EmbeddedTLB.scala 476:20]
      REG_3 <= 1'h0; // @[EmbeddedTLB.scala 476:28]
    end else begin
      REG_3 <= _GEN_5;
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_addr <= 39'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_addr <= io_in_req_bits_addr; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_size <= 3'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_size <= io_in_req_bits_size; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_cmd <= 4'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_cmd <= io_in_req_bits_cmd; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_wmask <= 8'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_wmask <= io_in_req_bits_wmask; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_req_wdata <= 64'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_req_wdata <= io_in_req_bits_wdata; // @[EmbeddedTLB.scala 608:31]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_hitVec <= 4'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_hitVec <= _T_214; // @[EmbeddedTLB.scala 610:34]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_miss <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_miss <= _T_219; // @[EmbeddedTLB.scala 611:32]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_hitWB <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_hitWB <= _T_286; // @[EmbeddedTLB.scala 612:33]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_loadPF <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_loadPF <= _T_318; // @[EmbeddedTLB.scala 613:34]
      end
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_1_storePF <= 1'h0; // @[EmbeddedTLB.scala 491:25]
      end else begin
        r_1_storePF <= _T_332; // @[EmbeddedTLB.scala 614:35]
      end
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_4 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush) begin // @[Pipeline.scala 27:20]
      REG_4 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_4 <= _GEN_19;
    end
    if (reset) begin // @[EmbeddedTLB.scala 505:22]
      state <= 1'h0; // @[EmbeddedTLB.scala 505:22]
    end else if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
      if (io_flush) begin // @[EmbeddedTLB.scala 520:19]
        state <= 1'h0; // @[EmbeddedTLB.scala 520:26]
      end
    end else if (_T_333) begin // @[EmbeddedTLB.scala 586:19]
      state <= _GEN_29;
    end else if (state) begin // @[EmbeddedTLB.scala 586:19]
      state <= _GEN_31;
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      r_2_addr <= out_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_2_size <= tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 495:16]
      end else begin
        r_2_size <= io_in_req_bits_size; // @[EmbeddedTLB.scala 576:18]
      end
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_2_cmd <= tlbExec_io_out_bits_cmd; // @[EmbeddedTLB.scala 495:16]
      end else begin
        r_2_cmd <= io_in_req_bits_cmd; // @[EmbeddedTLB.scala 576:18]
      end
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_2_wmask <= tlbExec_io_out_bits_wmask; // @[EmbeddedTLB.scala 495:16]
      end else begin
        r_2_wmask <= io_in_req_bits_wmask; // @[EmbeddedTLB.scala 576:18]
      end
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      if (~vmEnable) begin // @[EmbeddedTLB.scala 507:19]
        r_2_wdata <= tlbExec_io_out_bits_wdata; // @[EmbeddedTLB.scala 495:16]
      end else begin
        r_2_wdata <= io_in_req_bits_wdata; // @[EmbeddedTLB.scala 576:18]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  REG_2 = _RAND_2[38:0];
  _RAND_3 = {4{`RANDOM}};
  r__0 = _RAND_3[120:0];
  _RAND_4 = {4{`RANDOM}};
  r__1 = _RAND_4[120:0];
  _RAND_5 = {4{`RANDOM}};
  r__2 = _RAND_5[120:0];
  _RAND_6 = {4{`RANDOM}};
  r__3 = _RAND_6[120:0];
  _RAND_7 = {2{`RANDOM}};
  REG_5 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  REG_3 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_req_addr = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_req_size = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  r_1_req_cmd = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  r_1_req_wmask = _RAND_12[7:0];
  _RAND_13 = {2{`RANDOM}};
  r_1_req_wdata = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  r_1_hitVec = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  r_1_miss = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_hitWB = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_loadPF = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_1_storePF = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG_4 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  state = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  r_2_addr = _RAND_21[38:0];
  _RAND_22 = {1{`RANDOM}};
  r_2_size = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  r_2_cmd = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  r_2_wmask = _RAND_24[7:0];
  _RAND_25 = {2{`RANDOM}};
  r_2_wdata = _RAND_25[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_24 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_24) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 147:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 146:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 145:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 145:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 145:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 145:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 145:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module CacheStage2_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [18:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_dirty,
  output [18:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_dirty,
  output [18:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_dirty,
  output [18:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 176:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 176:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 176:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 178:64]
  reg  isForwardMetaReg; // @[Cache.scala 179:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 180:24 179:33 180:43]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 181:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 181:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 15:16 16:{19,23}]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 15:16 16:{19,23}]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 15:16 16:{19,23}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 185:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 187:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 187:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 187:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 187:61]
  wire [18:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[Cache.scala 189:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 192:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_39 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_42 = {_T_39,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 193:42]
  wire  _T_45 = ~metaWay_0_valid; // @[Cache.scala 195:45]
  wire  _T_46 = ~metaWay_1_valid; // @[Cache.scala 195:45]
  wire  _T_47 = ~metaWay_2_valid; // @[Cache.scala 195:45]
  wire  _T_48 = ~metaWay_3_valid; // @[Cache.scala 195:45]
  wire [3:0] invalidVec = {_T_48,_T_47,_T_46,_T_45}; // @[Cache.scala 195:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 196:34]
  wire [1:0] _T_52 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 199:8]
  wire [2:0] _T_53 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_52}; // @[Cache.scala 198:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_53}; // @[Cache.scala 197:33]
  wire [3:0] _T_54 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 202:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  wire [1:0] _T_59 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_61 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_63 = _T_59 + _T_61; // @[Bitwise.scala 47:55]
  wire  _T_65 = _T_63 > 3'h1; // @[Cache.scala 203:26]
  wire  _T_173 = io_in_bits_req_addr < 32'h40000000; // @[NutCore.scala 92:35]
  wire  _T_177 = io_in_bits_req_addr >= 32'h40600000 & io_in_bits_req_addr < 32'h41600000; // @[NutCore.scala 92:26]
  wire [9:0] _T_194 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_196 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_194; // @[Cache.scala 220:13]
  wire  isForwardData = io_in_valid & _T_196; // @[Cache.scala 219:35]
  reg  isForwardDataReg; // @[Cache.scala 222:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 223:24 222:33 223:43]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_203 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_203; // @[Cache.scala 231:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 230:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 229:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 229:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 229:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 229:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 229:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 215:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 213:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  assign io_out_bits_mmio = _T_173 | _T_177; // @[NutCore.scala 93:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 226:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 227:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 227:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 179:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 179:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 181:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 181:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_42;
    end
    if (reset) begin // @[Cache.scala 222:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 222:33]
    end else if (_T_12) begin // @[Cache.scala 224:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 224:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 16:23]
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:210 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 210:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fatal; // @[Cache.scala 210:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  REG = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage3_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [18:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_dirty,
  input  [18:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_dirty,
  input  [18:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_dirty,
  input  [18:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid,
  output [3:0]  io_cohResp_bits_cmd,
  output [63:0] io_cohResp_bits_rdata,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 257:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 257:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 257:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 257:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 257:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 257:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 258:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 258:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 258:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 258:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 258:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 258:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 261:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 261:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 262:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 263:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 264:26]
  wire  _T_6 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_6; // @[Cache.scala 265:39]
  wire  _T_7 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_7; // @[Cache.scala 266:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[Mux.scala 27:72]
  wire [18:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [18:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 277:49]
  wire [63:0] _T_50 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_51 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_52 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_53 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_54 = _T_50 | _T_51; // @[Mux.scala 27:72]
  wire [63:0] _T_55 = _T_54 | _T_52; // @[Mux.scala 27:72]
  wire [63:0] _T_56 = _T_55 | _T_53; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_56; // @[Cache.scala 279:21]
  wire [7:0] _T_69 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_77 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_79 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_81 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_83 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_84 = {_T_83,_T_81,_T_79,_T_77,_T_75,_T_73,_T_71,_T_69}; // @[Cat.scala 30:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_84 : 64'h0; // @[Cache.scala 280:21]
  reg [2:0] value; // @[Counter.scala 60:40]
  wire  _T_85 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_86 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 283:34]
  wire  _T_87 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_88 = io_in_bits_req_cmd == 4'h3 | _T_87; // @[Cache.scala 283:62]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_0 = _T_85 & (io_in_bits_req_cmd == 4'h3 | _T_87) ? _value_T_1 : value; // @[Cache.scala 283:85 Counter.scala 76:15 60:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 287:22]
  wire [63:0] _T_91 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_92 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_93 = dataRead & _T_92; // @[BitUtils.scala 32:36]
  wire [2:0] _T_98 = _T_88 ? value : addr_wordIndex; // @[Cache.scala 290:51]
  wire  metaHitWriteBus_req_valid = hitWrite & ~meta_dirty; // @[Cache.scala 293:22]
  reg [3:0] state; // @[Cache.scala 298:22]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 308:23]
  wire  _T_110 = state == 4'h3; // @[Cache.scala 310:39]
  wire  _T_111 = state == 4'h8; // @[Cache.scala 310:66]
  wire [2:0] _T_116 = _T_111 ? value_1 : value_2; // @[Cache.scala 311:33]
  wire  _T_118 = state2 == 2'h1; // @[Cache.scala 312:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_123 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_124 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_125 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_126 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_127 = _T_123 | _T_124; // @[Mux.scala 27:72]
  wire [63:0] _T_128 = _T_127 | _T_125; // @[Mux.scala 27:72]
  wire  _T_131 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_134 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_137 = hitReadBurst & io_out_ready; // @[Cache.scala 318:83]
  wire [1:0] _GEN_8 = _T_134 | io_cohResp_valid | hitReadBurst & io_out_ready ? 2'h0 : state2; // @[Cache.scala 318:{100,109} 308:23]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_140 = state == 4'h1; // @[Cache.scala 326:23]
  wire [2:0] _T_142 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 327:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_142; // @[Cache.scala 326:16]
  wire  _T_148 = state2 == 2'h2; // @[Cache.scala 333:89]
  reg  afterFirstRead; // @[Cache.scala 340:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_85 | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_154 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_156 = state == 4'h2; // @[Cache.scala 342:70]
  wire  readingFirst = ~afterFirstRead & _T_154 & state == 4'h2; // @[Cache.scala 342:60]
  wire  _T_159 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 344:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_160 = state == 4'h0; // @[Cache.scala 347:31]
  wire  _T_164 = _T_111 & _T_148; // @[Cache.scala 348:46]
  wire  _T_168 = _T_111 & io_cohResp_valid; // @[Cache.scala 350:49]
  reg [2:0] value_3; // @[Counter.scala 60:40]
  wire  wrap_wrap = value_3 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_1 = value_3 + 3'h1; // @[Counter.scala 76:24]
  wire  releaseLast = _T_168 & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire [2:0] _T_170 = releaseLast ? 3'h6 : 3'h0; // @[Cache.scala 351:54]
  wire [3:0] _T_171 = hit ? 4'hc : 4'h8; // @[Cache.scala 352:8]
  wire  respToL1Fire = _T_137 & _T_148; // @[Cache.scala 354:51]
  wire  _T_181 = (_T_160 | _T_164) & hitReadBurst & io_out_ready; // @[Cache.scala 355:112]
  reg [2:0] value_4; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = value_4 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_3 = value_4 + 3'h1; // @[Counter.scala 76:24]
  wire  respToL1Last = _T_181 & wrap_wrap_1; // @[Counter.scala 118:{17,24}]
  wire [3:0] _T_184 = hit ? 4'h8 : 4'h0; // @[Cache.scala 364:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[Cache.scala 369:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[Cache.scala 369:33]
  wire [3:0] _T_191 = meta_dirty ? 4'h3 : 4'h1; // @[Cache.scala 371:42]
  wire [3:0] _T_192 = mmio ? 4'h5 : _T_191; // @[Cache.scala 371:21]
  wire [3:0] _GEN_20 = miss | mmio ? _T_192 : state; // @[Cache.scala 370:49 371:15 298:22]
  wire  _T_194 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_196 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = _T_196 ? 4'h7 : state; // @[Cache.scala 298:22 376:{50,58}]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : value_1; // @[Cache.scala 379:48 Counter.scala 76:15 60:40]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[Cache.scala 298:22 380:{88,96}]
  wire [3:0] _GEN_29 = _T_134 ? 4'h2 : state; // @[Cache.scala 383:50 384:13 298:22]
  wire [2:0] _GEN_30 = _T_134 ? addr_wordIndex : value_1; // @[Cache.scala 383:50 385:25 Counter.scala 60:40]
  wire [2:0] _GEN_31 = _T_86 ? 3'h0 : _GEN_0; // @[Cache.scala 392:{52,75}]
  wire  _T_210 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_210 ? 4'h7 : state; // @[Cache.scala 298:22 393:{46,54}]
  wire  _GEN_33 = _T_154 | afterFirstRead; // @[Cache.scala 389:33 390:24 340:31]
  wire [2:0] _GEN_34 = _T_154 ? _value_T_7 : value_1; // @[Cache.scala 389:33 Counter.scala 76:15 60:40]
  wire [2:0] _GEN_35 = _T_154 ? _GEN_31 : _GEN_0; // @[Cache.scala 389:33]
  wire [3:0] _GEN_36 = _T_154 ? _GEN_32 : state; // @[Cache.scala 298:22 389:33]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_134 ? _value_T_11 : value_2; // @[Cache.scala 398:32 Counter.scala 76:15 60:40]
  wire  _T_213 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_213 & _T_134 ? 4'h4 : state; // @[Cache.scala 298:22 399:{65,73}]
  wire [3:0] _GEN_39 = _T_154 ? 4'h1 : state; // @[Cache.scala 298:22 402:{53,61}]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[Cache.scala 298:22 403:{76,84}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[Cache.scala 357:18 298:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[Cache.scala 357:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : value_2; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[Cache.scala 357:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : value_1; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [2:0] _GEN_47 = 4'h2 == state ? _GEN_35 : _GEN_0; // @[Cache.scala 357:18]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[Cache.scala 357:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? value_2 : _GEN_43; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[Cache.scala 357:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[Cache.scala 357:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_53 = 4'h1 == state ? _GEN_0 : _GEN_47; // @[Cache.scala 357:18]
  wire [2:0] _GEN_54 = 4'h1 == state ? value_2 : _GEN_49; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[Cache.scala 357:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? _GEN_28 : _GEN_50; // @[Cache.scala 357:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_58 = 4'h8 == state ? _GEN_0 : _GEN_53; // @[Cache.scala 357:18]
  wire [2:0] _GEN_59 = 4'h8 == state ? value_2 : _GEN_54; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [63:0] _T_222 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 406:67]
  wire [63:0] _T_223 = io_in_bits_req_wdata & _T_222; // @[BitUtils.scala 32:13]
  wire [63:0] _T_224 = ~_T_222; // @[BitUtils.scala 32:38]
  wire [63:0] _T_225 = io_mem_resp_bits_rdata & _T_224; // @[BitUtils.scala 32:36]
  wire  dataRefillWriteBus_req_valid = _T_156 & _T_154; // @[Cache.scala 408:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_210; // @[Cache.scala 416:61]
  wire  _T_247 = ~io_in_bits_req_cmd[0] & ~io_in_bits_req_cmd[3]; // @[SimpleBus.scala 73:26]
  wire [2:0] _T_249 = io_in_bits_req_cmd[0] ? 3'h5 : 3'h0; // @[Cache.scala 444:79]
  wire [2:0] _T_250 = _T_247 ? 3'h6 : _T_249; // @[Cache.scala 444:27]
  wire  _T_255 = state == 4'h7; // @[Cache.scala 450:48]
  wire  _T_274 = io_in_bits_req_cmd[0] | mmio ? _T_255 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 451:45]
  wire  _T_276 = probe ? 1'h0 : hit | _T_274; // @[Cache.scala 451:8]
  wire  _T_283 = miss ? _T_160 : _T_111 & releaseLast; // @[Cache.scala 458:53]
  wire  _T_292 = hit | io_in_bits_req_cmd[0] ? _T_85 : _T_255 & _GEN_12; // @[Cache.scala 459:8]
  Arbiter metaWriteArb ( // @[Cache.scala 257:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 258:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & (_T_160 & ~hitReadBurst) & ~miss & ~probe; // @[Cache.scala 462:79]
  assign io_out_valid = io_in_valid & _T_276; // @[Cache.scala 449:31]
  assign io_out_bits_cmd = {{1'd0}, _T_250}; // @[Cache.scala 444:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 443:29]
  assign io_isFinish = probe ? io_cohResp_valid & _T_283 : _T_292; // @[Cache.scala 458:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 310:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_116}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 413:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 423:23]
  assign io_mem_req_valid = _T_140 | _T_110 & state2 == 2'h2; // @[Cache.scala 333:48]
  assign io_mem_req_bits_addr = _T_140 ? raddr : waddr; // @[Cache.scala 328:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_128 | _T_126; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 332:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 338:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 336:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 336:20]
  assign io_mmio_req_bits_cmd = io_in_bits_req_cmd; // @[Cache.scala 336:20]
  assign io_mmio_req_bits_wmask = io_in_bits_req_wmask; // @[Cache.scala 336:20]
  assign io_mmio_req_bits_wdata = io_in_bits_req_wdata; // @[Cache.scala 336:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 337:22]
  assign io_cohResp_valid = state == 4'h0 & probe | _T_164; // @[Cache.scala 347:53]
  assign io_cohResp_bits_cmd = _T_111 ? {{1'd0}, _T_170} : _T_171; // @[Cache.scala 351:29]
  assign io_cohResp_bits_rdata = _T_128 | _T_126; // @[Mux.scala 27:72]
  assign io_dataReadRespToL1 = hitReadBurst & (_T_160 & io_out_ready | _T_164); // @[Cache.scala 463:39]
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[Cache.scala 293:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h1; // @[Cache.scala 294:16 97:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 292:29 SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_210; // @[Cache.scala 416:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 261:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 415:32 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 287:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_98}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = _T_91 | _T_93; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 288:29 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _T_156 & _T_154; // @[Cache.scala 408:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = _T_223 | _T_225; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 407:32 SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      value <= _GEN_0;
    end else if (4'h5 == state) begin // @[Cache.scala 357:18]
      value <= _GEN_0;
    end else if (4'h6 == state) begin // @[Cache.scala 357:18]
      value <= _GEN_0;
    end else begin
      value <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 298:22]
      state <= 4'h0; // @[Cache.scala 298:22]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      if (probe) begin // @[Cache.scala 362:20]
        if (io_cohResp_valid) begin // @[Cache.scala 363:34]
          state <= _T_184; // @[Cache.scala 364:17]
        end
      end else if (_T_137) begin // @[Cache.scala 367:50]
        state <= 4'h8; // @[Cache.scala 368:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (4'h5 == state) begin // @[Cache.scala 357:18]
      if (_T_194) begin // @[Cache.scala 375:48]
        state <= 4'h6; // @[Cache.scala 375:56]
      end
    end else if (4'h6 == state) begin // @[Cache.scala 357:18]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      if (probe) begin // @[Cache.scala 362:20]
        if (io_cohResp_valid) begin // @[Cache.scala 363:34]
          value_1 <= addr_wordIndex; // @[Cache.scala 365:29]
        end
      end else if (_T_137) begin // @[Cache.scala 367:50]
        value_1 <= _value_T_5; // @[Cache.scala 369:27]
      end
    end else if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
        value_1 <= _GEN_55;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 308:23]
      state2 <= 2'h0; // @[Cache.scala 308:23]
    end else if (2'h0 == state2) begin // @[Cache.scala 315:19]
      if (_T_131) begin // @[Cache.scala 316:53]
        state2 <= 2'h1; // @[Cache.scala 316:62]
      end
    end else if (2'h1 == state2) begin // @[Cache.scala 315:19]
      state2 <= 2'h2; // @[Cache.scala 317:35]
    end else if (2'h2 == state2) begin // @[Cache.scala 315:19]
      state2 <= _GEN_8;
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Cache.scala 340:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 340:31]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      afterFirstRead <= 1'h0; // @[Cache.scala 359:22]
    end else if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      alreadyOutFire <= 1'h0; // @[Cache.scala 360:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_159) begin // @[Reg.scala 16:19]
      if (mmio) begin // @[Cache.scala 343:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_3 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_168) begin // @[Counter.scala 118:17]
      value_3 <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_4 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_181) begin // @[Counter.scala 118:17]
      value_4 <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:268 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 268:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 268:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:465 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 465:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 465:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:466 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 466:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 466:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  value_3 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  value_4 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_9(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : io_in_1_bits_size; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_cmd = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_wmask = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  output        io_out_coh_req_ready,
  input         io_out_coh_req_valid,
  input  [31:0] io_out_coh_req_bits_addr,
  input  [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_valid,
  output [3:0]  io_out_coh_resp_bits_cmd,
  output [63:0] io_out_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 484:18]
  wire  s1_io_in_valid; // @[Cache.scala 484:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 484:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 484:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 484:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 484:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 484:18]
  wire  s1_io_out_ready; // @[Cache.scala 484:18]
  wire  s1_io_out_valid; // @[Cache.scala 484:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 484:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 484:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 484:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 484:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 484:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 484:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 484:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 484:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 484:18]
  wire  s2_clock; // @[Cache.scala 485:18]
  wire  s2_reset; // @[Cache.scala 485:18]
  wire  s2_io_in_ready; // @[Cache.scala 485:18]
  wire  s2_io_in_valid; // @[Cache.scala 485:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 485:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 485:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 485:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 485:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 485:18]
  wire  s2_io_out_ready; // @[Cache.scala 485:18]
  wire  s2_io_out_valid; // @[Cache.scala 485:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 485:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 485:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 485:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 485:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 485:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 485:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 485:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 485:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 485:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 485:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 485:18]
  wire  s3_clock; // @[Cache.scala 486:18]
  wire  s3_reset; // @[Cache.scala 486:18]
  wire  s3_io_in_ready; // @[Cache.scala 486:18]
  wire  s3_io_in_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 486:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 486:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 486:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 486:18]
  wire  s3_io_out_ready; // @[Cache.scala 486:18]
  wire  s3_io_out_valid; // @[Cache.scala 486:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_isFinish; // @[Cache.scala 486:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 486:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 486:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 486:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 486:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 486:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 486:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 486:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 486:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 486:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 486:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mmio_req_bits_cmd; // @[Cache.scala 486:18]
  wire [7:0] s3_io_mmio_req_bits_wmask; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mmio_req_bits_wdata; // @[Cache.scala 486:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 486:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 486:18]
  wire [3:0] s3_io_cohResp_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_cohResp_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 486:18]
  wire  metaArray_clock; // @[Cache.scala 487:25]
  wire  metaArray_reset; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 487:25]
  wire [6:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 487:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 487:25]
  wire [6:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 487:25]
  wire [18:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 487:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 487:25]
  wire  dataArray_clock; // @[Cache.scala 488:25]
  wire  dataArray_reset; // @[Cache.scala 488:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 488:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 488:25]
  wire [9:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 488:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 488:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 488:25]
  wire [9:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 488:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 488:25]
  wire [9:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 488:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 488:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 497:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 497:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 497:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 497:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 497:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 497:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 497:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 497:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 497:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 497:19]
  wire  arb_io_out_ready; // @[Cache.scala 497:19]
  wire  arb_io_out_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 497:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 497:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 497:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 497:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_req_size; // @[Reg.scala 15:16]
  reg [3:0] r_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_req_wdata; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_5 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_1_req_size; // @[Reg.scala 15:16]
  reg [3:0] r_1_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_1_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_1_req_wdata; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_0_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_0_dirty; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_1_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_1_dirty; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_2_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_2_dirty; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_3_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_3_data; // @[Reg.scala 15:16]
  reg  r_1_hit; // @[Reg.scala 15:16]
  reg [3:0] r_1_waymask; // @[Reg.scala 15:16]
  reg  r_1_mmio; // @[Reg.scala 15:16]
  reg  r_1_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] r_1_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] r_1_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_11 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  CacheStage1_1 s1 ( // @[Cache.scala 484:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2_1 s2 ( // @[Cache.scala 485:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3_1 s3 ( // @[Cache.scala 486:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(s3_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(s3_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(s3_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_cohResp_bits_cmd(s3_io_cohResp_bits_cmd),
    .io_cohResp_bits_rdata(s3_io_cohResp_bits_rdata),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 487:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 488:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 497:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 498:28]
  assign io_in_resp_valid = s3_io_out_valid & _T_11 ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 514:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 508:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 508:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 510:14]
  assign io_out_coh_req_ready = arb_io_in_0_ready; // @[Cache.scala 523:26]
  assign io_out_coh_resp_valid = s3_io_cohResp_valid; // @[Cache.scala 524:21]
  assign io_out_coh_resp_bits_cmd = s3_io_cohResp_bits_cmd; // @[Cache.scala 524:21]
  assign io_out_coh_resp_bits_rdata = s3_io_cohResp_bits_rdata; // @[Cache.scala 524:21]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_cmd = s3_io_mmio_req_bits_cmd; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_wmask = s3_io_mmio_req_bits_wmask; // @[Cache.scala 511:11]
  assign io_mmio_req_bits_wdata = s3_io_mmio_req_bits_wdata; // @[Cache.scala 511:11]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 500:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 500:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 500:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 500:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 500:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 500:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 532:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 533:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = r_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = r_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = r_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = r_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = r_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 539:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 542:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 541:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = r_1_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = r_1_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = r_1_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = r_1_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = r_1_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = r_1_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = r_1_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = r_1_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = r_1_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = r_1_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = r_1_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = r_1_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = r_1_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = r_1_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = r_1_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = r_1_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = r_1_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = r_1_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = r_1_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = r_1_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = r_1_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = r_1_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = r_1_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 508:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 534:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 510:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 511:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 511:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 511:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 532:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 532:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 536:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 533:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 533:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 534:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 534:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 537:18]
  assign arb_io_in_0_valid = io_out_coh_req_valid; // @[Cache.scala 522:24]
  assign arb_io_in_0_bits_addr = io_out_coh_req_bits_addr; // @[Cache.scala 519:19 SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_size = 3'h3; // @[Cache.scala 519:19 SimpleBus.scala 66:15]
  assign arb_io_in_0_bits_cmd = 4'h8; // @[Cache.scala 519:19 SimpleBus.scala 65:14]
  assign arb_io_in_0_bits_wmask = 8'hff; // @[Cache.scala 519:19 SimpleBus.scala 68:16]
  assign arb_io_in_0_bits_wdata = io_out_coh_req_bits_wdata; // @[Cache.scala 519:19 SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 498:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 500:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_size <= s1_io_out_bits_req_size; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_cmd <= s1_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wmask <= s1_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wdata <= s1_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_1 <= _GEN_9;
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_size <= s2_io_out_bits_req_size; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_cmd <= s2_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wmask <= s2_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wdata <= s2_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_hit <= s2_io_out_bits_hit; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  r_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  r_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  r_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  r_1_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  r_1_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  r_1_metas_0_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  r_1_metas_0_dirty = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_1_metas_1_tag = _RAND_14[18:0];
  _RAND_15 = {1{`RANDOM}};
  r_1_metas_1_dirty = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_metas_2_tag = _RAND_16[18:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_metas_2_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_1_metas_3_tag = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  r_1_metas_3_dirty = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  r_1_datas_0_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  r_1_datas_1_data = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  r_1_datas_2_data = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  r_1_datas_3_data = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  r_1_hit = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_1_waymask = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  r_1_mmio = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_1_isForwardData = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  r_1_forwardData_data_data = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  r_1_forwardData_waymask = _RAND_29[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready,
  output        io_imem_mem_req_valid,
  output [31:0] io_imem_mem_req_bits_addr,
  output [3:0]  io_imem_mem_req_bits_cmd,
  output [63:0] io_imem_mem_req_bits_wdata,
  input         io_imem_mem_resp_valid,
  input  [3:0]  io_imem_mem_resp_bits_cmd,
  input  [63:0] io_imem_mem_resp_bits_rdata,
  input         io_dmem_mem_req_ready,
  output        io_dmem_mem_req_valid,
  output [31:0] io_dmem_mem_req_bits_addr,
  output [3:0]  io_dmem_mem_req_bits_cmd,
  output [63:0] io_dmem_mem_req_bits_wdata,
  input         io_dmem_mem_resp_valid,
  input  [3:0]  io_dmem_mem_resp_bits_cmd,
  input  [63:0] io_dmem_mem_resp_bits_rdata,
  output        io_dmem_coh_req_ready,
  input         io_dmem_coh_req_valid,
  input  [31:0] io_dmem_coh_req_bits_addr,
  input  [63:0] io_dmem_coh_req_bits_wdata,
  output        io_dmem_coh_resp_valid,
  output [3:0]  io_dmem_coh_resp_bits_cmd,
  output [63:0] io_dmem_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [3:0]  io_mmio_resp_bits_cmd,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_frontend_req_ready,
  input         io_frontend_req_valid,
  input  [31:0] io_frontend_req_bits_addr,
  input  [2:0]  io_frontend_req_bits_size,
  input  [3:0]  io_frontend_req_bits_cmd,
  input  [7:0]  io_frontend_req_bits_wmask,
  input  [63:0] io_frontend_req_bits_wdata,
  input         io_frontend_resp_ready,
  output        io_frontend_resp_valid,
  output [3:0]  io_frontend_resp_bits_cmd,
  output [63:0] io_frontend_resp_bits_rdata,
  output [63:0] perfCnts_2,
  output [38:0] io_in_0_bits_decode_cf_pc,
  output [4:0]  io_wb_rfDest_0,
  input         io_extra_mtip,
  input         io_extra_meip_0,
  output        io_wb_rfWen_0,
  output [63:0] io_wb_WriteData_0,
  input         io_extra_msip,
  output        io_in_0_valid_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [63:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [63:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[NutCore.scala 106:24]
  wire  frontend_reset; // @[NutCore.scala 106:24]
  wire  frontend_io_imem_req_ready; // @[NutCore.scala 106:24]
  wire  frontend_io_imem_req_valid; // @[NutCore.scala 106:24]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[NutCore.scala 106:24]
  wire [86:0] frontend_io_imem_req_bits_user; // @[NutCore.scala 106:24]
  wire  frontend_io_imem_resp_ready; // @[NutCore.scala 106:24]
  wire  frontend_io_imem_resp_valid; // @[NutCore.scala 106:24]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[NutCore.scala 106:24]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_ready; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_valid; // @[NutCore.scala 106:24]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[NutCore.scala 106:24]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[NutCore.scala 106:24]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[NutCore.scala 106:24]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 106:24]
  wire [63:0] frontend_io_out_0_bits_cf_runahead_checkpoint_id; // @[NutCore.scala 106:24]
  wire [4:0] frontend_io_out_0_bits_cf_instrType; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[NutCore.scala 106:24]
  wire [3:0] frontend_io_out_0_bits_ctrl_fuType; // @[NutCore.scala 106:24]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[NutCore.scala 106:24]
  wire [2:0] frontend_io_out_0_bits_ctrl_funct3; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_ctrl_func24; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_ctrl_func23; // @[NutCore.scala 106:24]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[NutCore.scala 106:24]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[NutCore.scala 106:24]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc3; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[NutCore.scala 106:24]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[NutCore.scala 106:24]
  wire  frontend_io_out_0_bits_ctrl_isMou; // @[NutCore.scala 106:24]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[NutCore.scala 106:24]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[NutCore.scala 106:24]
  wire [3:0] frontend_io_flushVec; // @[NutCore.scala 106:24]
  wire [38:0] frontend_io_redirect_target; // @[NutCore.scala 106:24]
  wire  frontend_io_redirect_valid; // @[NutCore.scala 106:24]
  wire  frontend_io_ipf; // @[NutCore.scala 106:24]
  wire  frontend_flushICache; // @[NutCore.scala 106:24]
  wire  frontend_bpuUpdateReq_valid; // @[NutCore.scala 106:24]
  wire [38:0] frontend_bpuUpdateReq_pc; // @[NutCore.scala 106:24]
  wire  frontend_bpuUpdateReq_isMissPredict; // @[NutCore.scala 106:24]
  wire [38:0] frontend_bpuUpdateReq_actualTarget; // @[NutCore.scala 106:24]
  wire  frontend_bpuUpdateReq_actualTaken; // @[NutCore.scala 106:24]
  wire [6:0] frontend_bpuUpdateReq_fuOpType; // @[NutCore.scala 106:24]
  wire [1:0] frontend_bpuUpdateReq_btbType; // @[NutCore.scala 106:24]
  wire  frontend_bpuUpdateReq_isRVC; // @[NutCore.scala 106:24]
  wire  frontend_vmEnable; // @[NutCore.scala 106:24]
  wire [63:0] frontend_intrVec; // @[NutCore.scala 106:24]
  wire  frontend_flushTLB; // @[NutCore.scala 106:24]
  wire  backend_clock; // @[NutCore.scala 150:25]
  wire  backend_reset; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_ready; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_valid; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_in_0_bits_cf_instr; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_in_0_bits_cf_pc; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_in_0_bits_cf_pnpc; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_1; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_2; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_12; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_0; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_1; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_2; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_3; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_4; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_5; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_6; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_7; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_8; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_9; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_10; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_intrVec_11; // @[NutCore.scala 150:25]
  wire [3:0] backend_io_in_0_bits_cf_brIdx; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_in_0_bits_cf_runahead_checkpoint_id; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_0_bits_cf_instrType; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_ctrl_src1Type; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_ctrl_src2Type; // @[NutCore.scala 150:25]
  wire [3:0] backend_io_in_0_bits_ctrl_fuType; // @[NutCore.scala 150:25]
  wire [6:0] backend_io_in_0_bits_ctrl_fuOpType; // @[NutCore.scala 150:25]
  wire [2:0] backend_io_in_0_bits_ctrl_funct3; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_ctrl_func24; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_ctrl_func23; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc1; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc2; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc3; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_ctrl_rfWen; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfDest; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_bits_ctrl_isMou; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_in_0_bits_data_imm; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_ready; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_valid; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_in_1_bits_cf_instr; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_in_1_bits_cf_pc; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_in_1_bits_cf_pnpc; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_exceptionVec_1; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_exceptionVec_2; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_exceptionVec_12; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_0; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_1; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_2; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_3; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_4; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_5; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_6; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_7; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_8; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_9; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_10; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_intrVec_11; // @[NutCore.scala 150:25]
  wire [3:0] backend_io_in_1_bits_cf_brIdx; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_cf_crossPageIPFFix; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_in_1_bits_cf_runahead_checkpoint_id; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_1_bits_cf_instrType; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_ctrl_src1Type; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_ctrl_src2Type; // @[NutCore.scala 150:25]
  wire [3:0] backend_io_in_1_bits_ctrl_fuType; // @[NutCore.scala 150:25]
  wire [6:0] backend_io_in_1_bits_ctrl_fuOpType; // @[NutCore.scala 150:25]
  wire [2:0] backend_io_in_1_bits_ctrl_funct3; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_ctrl_func24; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_ctrl_func23; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_1_bits_ctrl_rfSrc1; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_1_bits_ctrl_rfSrc2; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_1_bits_ctrl_rfSrc3; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_ctrl_rfWen; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_in_1_bits_ctrl_rfDest; // @[NutCore.scala 150:25]
  wire  backend_io_in_1_bits_ctrl_isMou; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_in_1_bits_data_imm; // @[NutCore.scala 150:25]
  wire [1:0] backend_io_flush; // @[NutCore.scala 150:25]
  wire  backend_io_dmem_req_ready; // @[NutCore.scala 150:25]
  wire  backend_io_dmem_req_valid; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_dmem_req_bits_addr; // @[NutCore.scala 150:25]
  wire [2:0] backend_io_dmem_req_bits_size; // @[NutCore.scala 150:25]
  wire [3:0] backend_io_dmem_req_bits_cmd; // @[NutCore.scala 150:25]
  wire [7:0] backend_io_dmem_req_bits_wmask; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_dmem_req_bits_wdata; // @[NutCore.scala 150:25]
  wire  backend_io_dmem_resp_valid; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_dmem_resp_bits_rdata; // @[NutCore.scala 150:25]
  wire [1:0] backend_io_memMMU_imem_priviledgeMode; // @[NutCore.scala 150:25]
  wire [1:0] backend_io_memMMU_dmem_priviledgeMode; // @[NutCore.scala 150:25]
  wire  backend_io_memMMU_dmem_status_sum; // @[NutCore.scala 150:25]
  wire  backend_io_memMMU_dmem_status_mxr; // @[NutCore.scala 150:25]
  wire  backend_io_memMMU_dmem_loadPF; // @[NutCore.scala 150:25]
  wire  backend_io_memMMU_dmem_storePF; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_memMMU_dmem_addr; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_redirect_target; // @[NutCore.scala 150:25]
  wire  backend_io_redirect_valid; // @[NutCore.scala 150:25]
  wire  backend__T_408_0; // @[NutCore.scala 150:25]
  wire  backend_flushICache; // @[NutCore.scala 150:25]
  wire [63:0] backend_perfCnts_2; // @[NutCore.scala 150:25]
  wire [38:0] backend_io_in_0_bits_decode_cf_pc; // @[NutCore.scala 150:25]
  wire [63:0] backend_satp; // @[NutCore.scala 150:25]
  wire  backend_bpuUpdateReq_valid; // @[NutCore.scala 150:25]
  wire [38:0] backend_bpuUpdateReq_pc; // @[NutCore.scala 150:25]
  wire  backend_bpuUpdateReq_isMissPredict; // @[NutCore.scala 150:25]
  wire [38:0] backend_bpuUpdateReq_actualTarget; // @[NutCore.scala 150:25]
  wire  backend_bpuUpdateReq_actualTaken; // @[NutCore.scala 150:25]
  wire [6:0] backend_bpuUpdateReq_fuOpType; // @[NutCore.scala 150:25]
  wire [1:0] backend_bpuUpdateReq_btbType; // @[NutCore.scala 150:25]
  wire  backend_bpuUpdateReq_isRVC; // @[NutCore.scala 150:25]
  wire [4:0] backend_io_wb_rfDest_0; // @[NutCore.scala 150:25]
  wire  backend_ismmio; // @[NutCore.scala 150:25]
  wire  backend_io_extra_mtip; // @[NutCore.scala 150:25]
  wire  backend_amoReq; // @[NutCore.scala 150:25]
  wire  backend_io_extra_meip_0; // @[NutCore.scala 150:25]
  wire  backend_vmEnable; // @[NutCore.scala 150:25]
  wire  backend_io_wb_rfWen_0; // @[NutCore.scala 150:25]
  wire [63:0] backend_io_wb_WriteData_0; // @[NutCore.scala 150:25]
  wire [63:0] backend_intrVec; // @[NutCore.scala 150:25]
  wire  backend__T_407_0; // @[NutCore.scala 150:25]
  wire  backend_io_extra_msip; // @[NutCore.scala 150:25]
  wire  backend_flushTLB; // @[NutCore.scala 150:25]
  wire  backend_io_in_0_valid_0; // @[NutCore.scala 150:25]
  wire  mmioXbar_clock; // @[NutCore.scala 158:26]
  wire  mmioXbar_reset; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_in_0_req_ready; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_in_0_req_valid; // @[NutCore.scala 158:26]
  wire [31:0] mmioXbar_io_in_0_req_bits_addr; // @[NutCore.scala 158:26]
  wire [2:0] mmioXbar_io_in_0_req_bits_size; // @[NutCore.scala 158:26]
  wire [3:0] mmioXbar_io_in_0_req_bits_cmd; // @[NutCore.scala 158:26]
  wire [7:0] mmioXbar_io_in_0_req_bits_wmask; // @[NutCore.scala 158:26]
  wire [63:0] mmioXbar_io_in_0_req_bits_wdata; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_in_0_resp_valid; // @[NutCore.scala 158:26]
  wire [3:0] mmioXbar_io_in_0_resp_bits_cmd; // @[NutCore.scala 158:26]
  wire [63:0] mmioXbar_io_in_0_resp_bits_rdata; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_in_1_req_ready; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_in_1_req_valid; // @[NutCore.scala 158:26]
  wire [31:0] mmioXbar_io_in_1_req_bits_addr; // @[NutCore.scala 158:26]
  wire [2:0] mmioXbar_io_in_1_req_bits_size; // @[NutCore.scala 158:26]
  wire [3:0] mmioXbar_io_in_1_req_bits_cmd; // @[NutCore.scala 158:26]
  wire [7:0] mmioXbar_io_in_1_req_bits_wmask; // @[NutCore.scala 158:26]
  wire [63:0] mmioXbar_io_in_1_req_bits_wdata; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_in_1_resp_valid; // @[NutCore.scala 158:26]
  wire [3:0] mmioXbar_io_in_1_resp_bits_cmd; // @[NutCore.scala 158:26]
  wire [63:0] mmioXbar_io_in_1_resp_bits_rdata; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_out_req_ready; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_out_req_valid; // @[NutCore.scala 158:26]
  wire [31:0] mmioXbar_io_out_req_bits_addr; // @[NutCore.scala 158:26]
  wire [2:0] mmioXbar_io_out_req_bits_size; // @[NutCore.scala 158:26]
  wire [3:0] mmioXbar_io_out_req_bits_cmd; // @[NutCore.scala 158:26]
  wire [7:0] mmioXbar_io_out_req_bits_wmask; // @[NutCore.scala 158:26]
  wire [63:0] mmioXbar_io_out_req_bits_wdata; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_out_resp_ready; // @[NutCore.scala 158:26]
  wire  mmioXbar_io_out_resp_valid; // @[NutCore.scala 158:26]
  wire [3:0] mmioXbar_io_out_resp_bits_cmd; // @[NutCore.scala 158:26]
  wire [63:0] mmioXbar_io_out_resp_bits_rdata; // @[NutCore.scala 158:26]
  wire  dmemXbar_clock; // @[NutCore.scala 159:26]
  wire  dmemXbar_reset; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_0_req_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_0_req_valid; // @[NutCore.scala 159:26]
  wire [31:0] dmemXbar_io_in_0_req_bits_addr; // @[NutCore.scala 159:26]
  wire [2:0] dmemXbar_io_in_0_req_bits_size; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_in_0_req_bits_cmd; // @[NutCore.scala 159:26]
  wire [7:0] dmemXbar_io_in_0_req_bits_wmask; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_0_req_bits_wdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_0_resp_valid; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_0_resp_bits_rdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_1_req_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_1_req_valid; // @[NutCore.scala 159:26]
  wire [31:0] dmemXbar_io_in_1_req_bits_addr; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_in_1_req_bits_cmd; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_1_req_bits_wdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_1_resp_valid; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_1_resp_bits_rdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_2_req_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_2_req_valid; // @[NutCore.scala 159:26]
  wire [31:0] dmemXbar_io_in_2_req_bits_addr; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_in_2_req_bits_cmd; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_2_req_bits_wdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_2_resp_valid; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_2_resp_bits_rdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_3_req_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_3_req_valid; // @[NutCore.scala 159:26]
  wire [31:0] dmemXbar_io_in_3_req_bits_addr; // @[NutCore.scala 159:26]
  wire [2:0] dmemXbar_io_in_3_req_bits_size; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_in_3_req_bits_cmd; // @[NutCore.scala 159:26]
  wire [7:0] dmemXbar_io_in_3_req_bits_wmask; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_3_req_bits_wdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_3_resp_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_in_3_resp_valid; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_in_3_resp_bits_cmd; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_in_3_resp_bits_rdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_out_req_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_out_req_valid; // @[NutCore.scala 159:26]
  wire [31:0] dmemXbar_io_out_req_bits_addr; // @[NutCore.scala 159:26]
  wire [2:0] dmemXbar_io_out_req_bits_size; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_out_req_bits_cmd; // @[NutCore.scala 159:26]
  wire [7:0] dmemXbar_io_out_req_bits_wmask; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_out_req_bits_wdata; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_out_resp_ready; // @[NutCore.scala 159:26]
  wire  dmemXbar_io_out_resp_valid; // @[NutCore.scala 159:26]
  wire [3:0] dmemXbar_io_out_resp_bits_cmd; // @[NutCore.scala 159:26]
  wire [63:0] dmemXbar_io_out_resp_bits_rdata; // @[NutCore.scala 159:26]
  wire  itlb_clock; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_reset; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_in_req_ready; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_in_req_valid; // @[EmbeddedTLB.scala 425:13]
  wire [38:0] itlb_io_in_req_bits_addr; // @[EmbeddedTLB.scala 425:13]
  wire [86:0] itlb_io_in_req_bits_user; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_in_resp_ready; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_in_resp_valid; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] itlb_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 425:13]
  wire [86:0] itlb_io_in_resp_bits_user; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_out_req_ready; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_out_req_valid; // @[EmbeddedTLB.scala 425:13]
  wire [31:0] itlb_io_out_req_bits_addr; // @[EmbeddedTLB.scala 425:13]
  wire [2:0] itlb_io_out_req_bits_size; // @[EmbeddedTLB.scala 425:13]
  wire [86:0] itlb_io_out_req_bits_user; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_out_resp_ready; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_out_resp_valid; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] itlb_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 425:13]
  wire [86:0] itlb_io_out_resp_bits_user; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_mem_req_ready; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_mem_req_valid; // @[EmbeddedTLB.scala 425:13]
  wire [31:0] itlb_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 425:13]
  wire [3:0] itlb_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] itlb_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_mem_resp_valid; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] itlb_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_flush; // @[EmbeddedTLB.scala 425:13]
  wire [1:0] itlb_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_csrMMU_storePF; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_cacheEmpty; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_io_ipf; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] itlb_CSRSATP; // @[EmbeddedTLB.scala 425:13]
  wire  itlb_MOUFlushTLB; // @[EmbeddedTLB.scala 425:13]
  wire  Cache_clock; // @[Cache.scala 674:35]
  wire  Cache_reset; // @[Cache.scala 674:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 674:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 674:35]
  wire [2:0] Cache_io_in_req_bits_size; // @[Cache.scala 674:35]
  wire [86:0] Cache_io_in_req_bits_user; // @[Cache.scala 674:35]
  wire  Cache_io_in_resp_ready; // @[Cache.scala 674:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 674:35]
  wire [86:0] Cache_io_in_resp_bits_user; // @[Cache.scala 674:35]
  wire [1:0] Cache_io_flush; // @[Cache.scala 674:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 674:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 674:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 674:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  Cache_io_mmio_req_ready; // @[Cache.scala 674:35]
  wire  Cache_io_mmio_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_io_mmio_req_bits_addr; // @[Cache.scala 674:35]
  wire [2:0] Cache_io_mmio_req_bits_size; // @[Cache.scala 674:35]
  wire  Cache_io_mmio_resp_valid; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_mmio_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  Cache_io_empty; // @[Cache.scala 674:35]
  wire  Cache_MOUFlushICache; // @[Cache.scala 674:35]
  wire  dtlb_clock; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_reset; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_in_req_ready; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_in_req_valid; // @[EmbeddedTLB.scala 425:13]
  wire [38:0] dtlb_io_in_req_bits_addr; // @[EmbeddedTLB.scala 425:13]
  wire [2:0] dtlb_io_in_req_bits_size; // @[EmbeddedTLB.scala 425:13]
  wire [3:0] dtlb_io_in_req_bits_cmd; // @[EmbeddedTLB.scala 425:13]
  wire [7:0] dtlb_io_in_req_bits_wmask; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_io_in_req_bits_wdata; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_in_resp_valid; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_out_req_ready; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_out_req_valid; // @[EmbeddedTLB.scala 425:13]
  wire [31:0] dtlb_io_out_req_bits_addr; // @[EmbeddedTLB.scala 425:13]
  wire [2:0] dtlb_io_out_req_bits_size; // @[EmbeddedTLB.scala 425:13]
  wire [3:0] dtlb_io_out_req_bits_cmd; // @[EmbeddedTLB.scala 425:13]
  wire [7:0] dtlb_io_out_req_bits_wmask; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_io_out_req_bits_wdata; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_out_resp_valid; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_mem_req_ready; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_mem_req_valid; // @[EmbeddedTLB.scala 425:13]
  wire [31:0] dtlb_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 425:13]
  wire [3:0] dtlb_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_mem_resp_valid; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_flush; // @[EmbeddedTLB.scala 425:13]
  wire [1:0] dtlb_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_csrMMU_status_sum; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_io_csrMMU_storePF; // @[EmbeddedTLB.scala 425:13]
  wire [38:0] dtlb_io_csrMMU_addr; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb__T_408_0; // @[EmbeddedTLB.scala 425:13]
  wire [63:0] dtlb_CSRSATP; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_ismmio_0; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_ISAMO; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_vmEnable_0; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb__T_407_0; // @[EmbeddedTLB.scala 425:13]
  wire  dtlb_MOUFlushTLB; // @[EmbeddedTLB.scala 425:13]
  wire  Cache_1_clock; // @[Cache.scala 674:35]
  wire  Cache_1_reset; // @[Cache.scala 674:35]
  wire  Cache_1_io_in_req_ready; // @[Cache.scala 674:35]
  wire  Cache_1_io_in_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_1_io_in_req_bits_addr; // @[Cache.scala 674:35]
  wire [2:0] Cache_1_io_in_req_bits_size; // @[Cache.scala 674:35]
  wire [3:0] Cache_1_io_in_req_bits_cmd; // @[Cache.scala 674:35]
  wire [7:0] Cache_1_io_in_req_bits_wmask; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_in_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_in_resp_ready; // @[Cache.scala 674:35]
  wire  Cache_1_io_in_resp_valid; // @[Cache.scala 674:35]
  wire [3:0] Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_out_mem_req_ready; // @[Cache.scala 674:35]
  wire  Cache_1_io_out_mem_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_1_io_out_mem_req_bits_addr; // @[Cache.scala 674:35]
  wire [3:0] Cache_1_io_out_mem_req_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_out_mem_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_out_mem_resp_valid; // @[Cache.scala 674:35]
  wire [3:0] Cache_1_io_out_mem_resp_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_out_mem_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_out_coh_req_ready; // @[Cache.scala 674:35]
  wire  Cache_1_io_out_coh_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_1_io_out_coh_req_bits_addr; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_out_coh_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_out_coh_resp_valid; // @[Cache.scala 674:35]
  wire [3:0] Cache_1_io_out_coh_resp_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_out_coh_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_mmio_req_ready; // @[Cache.scala 674:35]
  wire  Cache_1_io_mmio_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 674:35]
  wire [2:0] Cache_1_io_mmio_req_bits_size; // @[Cache.scala 674:35]
  wire [3:0] Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 674:35]
  wire [7:0] Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_1_io_mmio_resp_valid; // @[Cache.scala 674:35]
  wire [63:0] Cache_1_io_mmio_resp_bits_rdata; // @[Cache.scala 674:35]
  reg [63:0] REG__0_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__0_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__0_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__0_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__0_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__0_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__1_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__1_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__1_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__1_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__2_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__2_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__2_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__2_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__3_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__3_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__3_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__3_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__4_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__4_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__4_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__4_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__4_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__4_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__4_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__4_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__4_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__4_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__4_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__4_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__4_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__4_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__4_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__4_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__4_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__4_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__4_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__4_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__4_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__5_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__5_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__5_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__5_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__5_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__5_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__5_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__5_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__5_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__5_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__5_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__5_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__5_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__5_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__5_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__5_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__5_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__5_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__5_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__5_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__5_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__6_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__6_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__6_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__6_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__6_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__6_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__6_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__6_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__6_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__6_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__6_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__6_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__6_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__6_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__6_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__6_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__6_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__6_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__6_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__6_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__6_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__7_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__7_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__7_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__7_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__7_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__7_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__7_cf_instrType; // @[PipelineVector.scala 29:29]
  reg  REG__7_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__7_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__7_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__7_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__7_ctrl_funct3; // @[PipelineVector.scala 29:29]
  reg  REG__7_ctrl_func24; // @[PipelineVector.scala 29:29]
  reg  REG__7_ctrl_func23; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__7_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__7_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__7_ctrl_rfSrc3; // @[PipelineVector.scala 29:29]
  reg  REG__7_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__7_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  REG__7_ctrl_isMou; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__7_data_imm; // @[PipelineVector.scala 29:29]
  reg [2:0] REG_1; // @[PipelineVector.scala 30:33]
  reg [2:0] REG_2; // @[PipelineVector.scala 31:33]
  wire [2:0] _T_3 = REG_1 + 3'h1; // @[PipelineVector.scala 33:63]
  wire [2:0] _T_6 = REG_1 + 3'h2; // @[PipelineVector.scala 33:63]
  wire  _T_9 = _T_3 != REG_2 & _T_6 != REG_2; // @[PipelineVector.scala 33:124]
  wire  _WIRE_9_0 = frontend_io_out_0_valid; // @[PipelineVector.scala 36:27 37:20]
  wire [1:0] _T_10 = {{1'd0}, _WIRE_9_0}; // @[PipelineVector.scala 40:46]
  wire  _T_11 = _T_10 >= 2'h1; // @[PipelineVector.scala 41:53]
  wire  _T_12 = _T_10 >= 2'h2; // @[PipelineVector.scala 41:53]
  wire  _T_13 = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_16 = {{1'd0}, REG_1}; // @[PipelineVector.scala 45:45]
  wire [63:0] _T_18_cf_instr = _WIRE_9_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_18_cf_pc = _WIRE_9_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_18_cf_pnpc = _WIRE_9_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_0 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_0 : frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_1 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_1 : frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_2 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_2 : frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_3 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_3 : frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_4 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_4 : frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_5 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_5 : frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_6 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_6 : frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_7 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_7 : frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_8 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_8 : frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_9 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_9 : frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_10 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_10 : frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_11 = _WIRE_9_0 ? frontend_io_out_0_bits_cf_intrVec_11 : frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_18_cf_brIdx = _WIRE_9_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_18_cf_runahead_checkpoint_id = _WIRE_9_0 ? frontend_io_out_0_bits_cf_runahead_checkpoint_id : 64'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_cf_instrType = _WIRE_9_0 ? frontend_io_out_0_bits_cf_instrType : 5'h0; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_src1Type = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_src1Type : 1'h1; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_src2Type = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_src2Type : 1'h1; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_18_ctrl_fuType = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_fuType : 4'h1; // @[PipelineVector.scala 45:69]
  wire [6:0] _T_18_ctrl_fuOpType = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[PipelineVector.scala 45:69]
  wire [2:0] _T_18_ctrl_funct3 = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_funct3 : 3'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc1 = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc2 = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc3 = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_rfSrc3 : 5'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfDest = _WIRE_9_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_18_data_imm = _WIRE_9_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[PipelineVector.scala 45:69]
  wire [63:0] _GEN_24 = 3'h0 == _T_16[2:0] ? _T_18_data_imm : REG__0_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_25 = 3'h1 == _T_16[2:0] ? _T_18_data_imm : REG__1_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_26 = 3'h2 == _T_16[2:0] ? _T_18_data_imm : REG__2_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_27 = 3'h3 == _T_16[2:0] ? _T_18_data_imm : REG__3_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_28 = 3'h4 == _T_16[2:0] ? _T_18_data_imm : REG__4_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_29 = 3'h5 == _T_16[2:0] ? _T_18_data_imm : REG__5_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_30 = 3'h6 == _T_16[2:0] ? _T_18_data_imm : REG__6_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_31 = 3'h7 == _T_16[2:0] ? _T_18_data_imm : REG__7_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_56 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__0_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_57 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__1_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_58 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__2_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_59 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__3_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_60 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__4_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_61 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__5_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_62 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__6_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_63 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_isMou : REG__7_ctrl_isMou; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_112 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_113 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_114 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_115 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_116 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__4_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_117 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__5_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_118 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__6_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_119 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_rfDest : REG__7_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_120 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_121 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_122 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_123 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_124 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__4_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_125 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__5_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_126 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__6_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_127 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_rfWen : REG__7_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_128 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__0_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_129 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__1_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_130 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__2_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_131 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__3_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_132 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__4_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_133 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__5_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_134 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__6_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_135 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_rfSrc3 : REG__7_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_136 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_137 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_138 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_139 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_140 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__4_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_141 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__5_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_142 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__6_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_143 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_rfSrc2 : REG__7_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_144 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_145 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_146 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_147 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_148 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__4_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_149 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__5_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_150 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__6_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_151 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_rfSrc1 : REG__7_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_152 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__0_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_153 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__1_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_154 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__2_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_155 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__3_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_156 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__4_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_157 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__5_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_158 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__6_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_159 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func23 : REG__7_ctrl_func23; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_160 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__0_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_161 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__1_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_162 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__2_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_163 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__3_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_164 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__4_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_165 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__5_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_166 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__6_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_167 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_ctrl_func24 : REG__7_ctrl_func24; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_168 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__0_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_169 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__1_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_170 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__2_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_171 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__3_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_172 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__4_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_173 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__5_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_174 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__6_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_175 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_funct3 : REG__7_ctrl_funct3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_176 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_177 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_178 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_179 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_180 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__4_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_181 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__5_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_182 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__6_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_183 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_fuOpType : REG__7_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_184 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_185 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_186 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_187 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_188 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__4_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_189 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__5_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_190 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__6_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_191 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_fuType : REG__7_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_192 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_193 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_194 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_195 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_196 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__4_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_197 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__5_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_198 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__6_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_199 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_src2Type : REG__7_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_200 = 3'h0 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_201 = 3'h1 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_202 = 3'h2 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_203 = 3'h3 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_204 = 3'h4 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__4_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_205 = 3'h5 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__5_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_206 = 3'h6 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__6_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_207 = 3'h7 == _T_16[2:0] ? _T_18_ctrl_src1Type : REG__7_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_208 = 3'h0 == _T_16[2:0] ? _T_18_cf_instrType : REG__0_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_209 = 3'h1 == _T_16[2:0] ? _T_18_cf_instrType : REG__1_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_210 = 3'h2 == _T_16[2:0] ? _T_18_cf_instrType : REG__2_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_211 = 3'h3 == _T_16[2:0] ? _T_18_cf_instrType : REG__3_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_212 = 3'h4 == _T_16[2:0] ? _T_18_cf_instrType : REG__4_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_213 = 3'h5 == _T_16[2:0] ? _T_18_cf_instrType : REG__5_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_214 = 3'h6 == _T_16[2:0] ? _T_18_cf_instrType : REG__6_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_215 = 3'h7 == _T_16[2:0] ? _T_18_cf_instrType : REG__7_cf_instrType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_224 = 3'h0 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_225 = 3'h1 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__1_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_226 = 3'h2 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__2_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_227 = 3'h3 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__3_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_228 = 3'h4 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__4_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_229 = 3'h5 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__5_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_230 = 3'h6 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__6_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_231 = 3'h7 == _T_16[2:0] ? _T_18_cf_runahead_checkpoint_id : REG__7_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_232 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_233 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_234 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_235 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_236 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__4_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_237 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__5_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_238 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__6_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_239 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    REG__7_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_248 = 3'h0 == _T_16[2:0] ? _T_18_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_249 = 3'h1 == _T_16[2:0] ? _T_18_cf_brIdx : REG__1_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_250 = 3'h2 == _T_16[2:0] ? _T_18_cf_brIdx : REG__2_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_251 = 3'h3 == _T_16[2:0] ? _T_18_cf_brIdx : REG__3_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_252 = 3'h4 == _T_16[2:0] ? _T_18_cf_brIdx : REG__4_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_253 = 3'h5 == _T_16[2:0] ? _T_18_cf_brIdx : REG__5_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_254 = 3'h6 == _T_16[2:0] ? _T_18_cf_brIdx : REG__6_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_255 = 3'h7 == _T_16[2:0] ? _T_18_cf_brIdx : REG__7_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_256 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_257 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_258 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_259 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_260 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__4_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_261 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__5_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_262 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__6_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_263 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_0 : REG__7_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_264 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_265 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_266 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_267 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_268 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__4_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_269 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__5_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_270 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__6_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_271 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_1 : REG__7_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_272 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_273 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_274 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_275 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_276 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__4_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_277 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__5_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_278 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__6_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_279 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_2 : REG__7_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_280 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_281 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_282 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_283 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_284 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__4_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_285 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__5_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_286 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__6_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_287 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_3 : REG__7_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_288 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_289 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_290 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_291 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_292 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__4_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_293 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__5_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_294 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__6_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_295 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_4 : REG__7_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_296 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_297 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_298 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_299 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_300 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__4_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_301 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__5_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_302 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__6_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_303 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_5 : REG__7_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_304 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_305 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_306 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_307 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_308 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__4_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_309 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__5_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_310 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__6_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_311 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_6 : REG__7_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_312 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_313 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_314 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_315 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_316 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__4_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_317 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__5_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_318 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__6_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_319 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_7 : REG__7_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_320 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_321 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_322 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_323 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_324 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__4_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_325 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__5_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_326 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__6_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_327 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_8 : REG__7_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_328 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_329 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_330 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_331 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_332 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__4_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_333 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__5_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_334 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__6_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_335 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_9 : REG__7_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_336 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_337 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_338 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_339 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_340 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__4_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_341 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__5_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_342 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__6_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_343 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_10 : REG__7_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_344 = 3'h0 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_345 = 3'h1 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_346 = 3'h2 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_347 = 3'h3 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_348 = 3'h4 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__4_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_349 = 3'h5 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__5_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_350 = 3'h6 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__6_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_351 = 3'h7 == _T_16[2:0] ? _T_18_cf_intrVec_11 : REG__7_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_360 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_361 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_362 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_363 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_364 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__4_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_365 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__5_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_366 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__6_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_367 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_1 : REG__7_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_368 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_369 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_370 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_371 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_372 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__4_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_373 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__5_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_374 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__6_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_375 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_2 : REG__7_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_448 = 3'h0 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_449 = 3'h1 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_450 = 3'h2 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_451 = 3'h3 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_452 = 3'h4 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__4_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_453 = 3'h5 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__5_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_454 = 3'h6 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__6_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_455 = 3'h7 == _T_16[2:0] ? _WIRE_9_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    REG__7_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_504 = 3'h0 == _T_16[2:0] ? _T_18_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_505 = 3'h1 == _T_16[2:0] ? _T_18_cf_pnpc : REG__1_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_506 = 3'h2 == _T_16[2:0] ? _T_18_cf_pnpc : REG__2_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_507 = 3'h3 == _T_16[2:0] ? _T_18_cf_pnpc : REG__3_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_508 = 3'h4 == _T_16[2:0] ? _T_18_cf_pnpc : REG__4_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_509 = 3'h5 == _T_16[2:0] ? _T_18_cf_pnpc : REG__5_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_510 = 3'h6 == _T_16[2:0] ? _T_18_cf_pnpc : REG__6_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_511 = 3'h7 == _T_16[2:0] ? _T_18_cf_pnpc : REG__7_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_512 = 3'h0 == _T_16[2:0] ? _T_18_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_513 = 3'h1 == _T_16[2:0] ? _T_18_cf_pc : REG__1_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_514 = 3'h2 == _T_16[2:0] ? _T_18_cf_pc : REG__2_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_515 = 3'h3 == _T_16[2:0] ? _T_18_cf_pc : REG__3_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_516 = 3'h4 == _T_16[2:0] ? _T_18_cf_pc : REG__4_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_517 = 3'h5 == _T_16[2:0] ? _T_18_cf_pc : REG__5_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_518 = 3'h6 == _T_16[2:0] ? _T_18_cf_pc : REG__6_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_519 = 3'h7 == _T_16[2:0] ? _T_18_cf_pc : REG__7_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_520 = 3'h0 == _T_16[2:0] ? _T_18_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_521 = 3'h1 == _T_16[2:0] ? _T_18_cf_instr : REG__1_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_522 = 3'h2 == _T_16[2:0] ? _T_18_cf_instr : REG__2_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_523 = 3'h3 == _T_16[2:0] ? _T_18_cf_instr : REG__3_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_524 = 3'h4 == _T_16[2:0] ? _T_18_cf_instr : REG__4_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_525 = 3'h5 == _T_16[2:0] ? _T_18_cf_instr : REG__5_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_526 = 3'h6 == _T_16[2:0] ? _T_18_cf_instr : REG__6_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_527 = 3'h7 == _T_16[2:0] ? _T_18_cf_instr : REG__7_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_552 = _T_11 ? _GEN_24 : REG__0_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_553 = _T_11 ? _GEN_25 : REG__1_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_554 = _T_11 ? _GEN_26 : REG__2_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_555 = _T_11 ? _GEN_27 : REG__3_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_556 = _T_11 ? _GEN_28 : REG__4_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_557 = _T_11 ? _GEN_29 : REG__5_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_558 = _T_11 ? _GEN_30 : REG__6_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_559 = _T_11 ? _GEN_31 : REG__7_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_584 = _T_11 ? _GEN_56 : REG__0_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_585 = _T_11 ? _GEN_57 : REG__1_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_586 = _T_11 ? _GEN_58 : REG__2_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_587 = _T_11 ? _GEN_59 : REG__3_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_588 = _T_11 ? _GEN_60 : REG__4_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_589 = _T_11 ? _GEN_61 : REG__5_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_590 = _T_11 ? _GEN_62 : REG__6_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_591 = _T_11 ? _GEN_63 : REG__7_ctrl_isMou; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_640 = _T_11 ? _GEN_112 : REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_641 = _T_11 ? _GEN_113 : REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_642 = _T_11 ? _GEN_114 : REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_643 = _T_11 ? _GEN_115 : REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_644 = _T_11 ? _GEN_116 : REG__4_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_645 = _T_11 ? _GEN_117 : REG__5_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_646 = _T_11 ? _GEN_118 : REG__6_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_647 = _T_11 ? _GEN_119 : REG__7_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_648 = _T_11 ? _GEN_120 : REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_649 = _T_11 ? _GEN_121 : REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_650 = _T_11 ? _GEN_122 : REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_651 = _T_11 ? _GEN_123 : REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_652 = _T_11 ? _GEN_124 : REG__4_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_653 = _T_11 ? _GEN_125 : REG__5_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_654 = _T_11 ? _GEN_126 : REG__6_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_655 = _T_11 ? _GEN_127 : REG__7_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_656 = _T_11 ? _GEN_128 : REG__0_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_657 = _T_11 ? _GEN_129 : REG__1_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_658 = _T_11 ? _GEN_130 : REG__2_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_659 = _T_11 ? _GEN_131 : REG__3_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_660 = _T_11 ? _GEN_132 : REG__4_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_661 = _T_11 ? _GEN_133 : REG__5_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_662 = _T_11 ? _GEN_134 : REG__6_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_663 = _T_11 ? _GEN_135 : REG__7_ctrl_rfSrc3; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_664 = _T_11 ? _GEN_136 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_665 = _T_11 ? _GEN_137 : REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_666 = _T_11 ? _GEN_138 : REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_667 = _T_11 ? _GEN_139 : REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_668 = _T_11 ? _GEN_140 : REG__4_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_669 = _T_11 ? _GEN_141 : REG__5_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_670 = _T_11 ? _GEN_142 : REG__6_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_671 = _T_11 ? _GEN_143 : REG__7_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_672 = _T_11 ? _GEN_144 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_673 = _T_11 ? _GEN_145 : REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_674 = _T_11 ? _GEN_146 : REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_675 = _T_11 ? _GEN_147 : REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_676 = _T_11 ? _GEN_148 : REG__4_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_677 = _T_11 ? _GEN_149 : REG__5_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_678 = _T_11 ? _GEN_150 : REG__6_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_679 = _T_11 ? _GEN_151 : REG__7_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_680 = _T_11 ? _GEN_152 : REG__0_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_681 = _T_11 ? _GEN_153 : REG__1_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_682 = _T_11 ? _GEN_154 : REG__2_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_683 = _T_11 ? _GEN_155 : REG__3_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_684 = _T_11 ? _GEN_156 : REG__4_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_685 = _T_11 ? _GEN_157 : REG__5_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_686 = _T_11 ? _GEN_158 : REG__6_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_687 = _T_11 ? _GEN_159 : REG__7_ctrl_func23; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_688 = _T_11 ? _GEN_160 : REG__0_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_689 = _T_11 ? _GEN_161 : REG__1_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_690 = _T_11 ? _GEN_162 : REG__2_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_691 = _T_11 ? _GEN_163 : REG__3_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_692 = _T_11 ? _GEN_164 : REG__4_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_693 = _T_11 ? _GEN_165 : REG__5_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_694 = _T_11 ? _GEN_166 : REG__6_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_695 = _T_11 ? _GEN_167 : REG__7_ctrl_func24; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_696 = _T_11 ? _GEN_168 : REG__0_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_697 = _T_11 ? _GEN_169 : REG__1_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_698 = _T_11 ? _GEN_170 : REG__2_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_699 = _T_11 ? _GEN_171 : REG__3_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_700 = _T_11 ? _GEN_172 : REG__4_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_701 = _T_11 ? _GEN_173 : REG__5_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_702 = _T_11 ? _GEN_174 : REG__6_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_703 = _T_11 ? _GEN_175 : REG__7_ctrl_funct3; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_704 = _T_11 ? _GEN_176 : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_705 = _T_11 ? _GEN_177 : REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_706 = _T_11 ? _GEN_178 : REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_707 = _T_11 ? _GEN_179 : REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_708 = _T_11 ? _GEN_180 : REG__4_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_709 = _T_11 ? _GEN_181 : REG__5_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_710 = _T_11 ? _GEN_182 : REG__6_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_711 = _T_11 ? _GEN_183 : REG__7_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_712 = _T_11 ? _GEN_184 : REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_713 = _T_11 ? _GEN_185 : REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_714 = _T_11 ? _GEN_186 : REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_715 = _T_11 ? _GEN_187 : REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_716 = _T_11 ? _GEN_188 : REG__4_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_717 = _T_11 ? _GEN_189 : REG__5_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_718 = _T_11 ? _GEN_190 : REG__6_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_719 = _T_11 ? _GEN_191 : REG__7_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_720 = _T_11 ? _GEN_192 : REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_721 = _T_11 ? _GEN_193 : REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_722 = _T_11 ? _GEN_194 : REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_723 = _T_11 ? _GEN_195 : REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_724 = _T_11 ? _GEN_196 : REG__4_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_725 = _T_11 ? _GEN_197 : REG__5_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_726 = _T_11 ? _GEN_198 : REG__6_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_727 = _T_11 ? _GEN_199 : REG__7_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_728 = _T_11 ? _GEN_200 : REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_729 = _T_11 ? _GEN_201 : REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_730 = _T_11 ? _GEN_202 : REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_731 = _T_11 ? _GEN_203 : REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_732 = _T_11 ? _GEN_204 : REG__4_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_733 = _T_11 ? _GEN_205 : REG__5_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_734 = _T_11 ? _GEN_206 : REG__6_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_735 = _T_11 ? _GEN_207 : REG__7_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_736 = _T_11 ? _GEN_208 : REG__0_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_737 = _T_11 ? _GEN_209 : REG__1_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_738 = _T_11 ? _GEN_210 : REG__2_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_739 = _T_11 ? _GEN_211 : REG__3_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_740 = _T_11 ? _GEN_212 : REG__4_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_741 = _T_11 ? _GEN_213 : REG__5_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_742 = _T_11 ? _GEN_214 : REG__6_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_743 = _T_11 ? _GEN_215 : REG__7_cf_instrType; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_752 = _T_11 ? _GEN_224 : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_753 = _T_11 ? _GEN_225 : REG__1_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_754 = _T_11 ? _GEN_226 : REG__2_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_755 = _T_11 ? _GEN_227 : REG__3_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_756 = _T_11 ? _GEN_228 : REG__4_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_757 = _T_11 ? _GEN_229 : REG__5_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_758 = _T_11 ? _GEN_230 : REG__6_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_759 = _T_11 ? _GEN_231 : REG__7_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_760 = _T_11 ? _GEN_232 : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_761 = _T_11 ? _GEN_233 : REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_762 = _T_11 ? _GEN_234 : REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_763 = _T_11 ? _GEN_235 : REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_764 = _T_11 ? _GEN_236 : REG__4_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_765 = _T_11 ? _GEN_237 : REG__5_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_766 = _T_11 ? _GEN_238 : REG__6_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_767 = _T_11 ? _GEN_239 : REG__7_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_776 = _T_11 ? _GEN_248 : REG__0_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_777 = _T_11 ? _GEN_249 : REG__1_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_778 = _T_11 ? _GEN_250 : REG__2_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_779 = _T_11 ? _GEN_251 : REG__3_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_780 = _T_11 ? _GEN_252 : REG__4_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_781 = _T_11 ? _GEN_253 : REG__5_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_782 = _T_11 ? _GEN_254 : REG__6_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_783 = _T_11 ? _GEN_255 : REG__7_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_784 = _T_11 ? _GEN_256 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_785 = _T_11 ? _GEN_257 : REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_786 = _T_11 ? _GEN_258 : REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_787 = _T_11 ? _GEN_259 : REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_788 = _T_11 ? _GEN_260 : REG__4_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_789 = _T_11 ? _GEN_261 : REG__5_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_790 = _T_11 ? _GEN_262 : REG__6_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_791 = _T_11 ? _GEN_263 : REG__7_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_792 = _T_11 ? _GEN_264 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_793 = _T_11 ? _GEN_265 : REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_794 = _T_11 ? _GEN_266 : REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_795 = _T_11 ? _GEN_267 : REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_796 = _T_11 ? _GEN_268 : REG__4_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_797 = _T_11 ? _GEN_269 : REG__5_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_798 = _T_11 ? _GEN_270 : REG__6_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_799 = _T_11 ? _GEN_271 : REG__7_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_800 = _T_11 ? _GEN_272 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_801 = _T_11 ? _GEN_273 : REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_802 = _T_11 ? _GEN_274 : REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_803 = _T_11 ? _GEN_275 : REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_804 = _T_11 ? _GEN_276 : REG__4_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_805 = _T_11 ? _GEN_277 : REG__5_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_806 = _T_11 ? _GEN_278 : REG__6_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_807 = _T_11 ? _GEN_279 : REG__7_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_808 = _T_11 ? _GEN_280 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_809 = _T_11 ? _GEN_281 : REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_810 = _T_11 ? _GEN_282 : REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_811 = _T_11 ? _GEN_283 : REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_812 = _T_11 ? _GEN_284 : REG__4_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_813 = _T_11 ? _GEN_285 : REG__5_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_814 = _T_11 ? _GEN_286 : REG__6_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_815 = _T_11 ? _GEN_287 : REG__7_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_816 = _T_11 ? _GEN_288 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_817 = _T_11 ? _GEN_289 : REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_818 = _T_11 ? _GEN_290 : REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_819 = _T_11 ? _GEN_291 : REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_820 = _T_11 ? _GEN_292 : REG__4_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_821 = _T_11 ? _GEN_293 : REG__5_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_822 = _T_11 ? _GEN_294 : REG__6_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_823 = _T_11 ? _GEN_295 : REG__7_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_824 = _T_11 ? _GEN_296 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_825 = _T_11 ? _GEN_297 : REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_826 = _T_11 ? _GEN_298 : REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_827 = _T_11 ? _GEN_299 : REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_828 = _T_11 ? _GEN_300 : REG__4_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_829 = _T_11 ? _GEN_301 : REG__5_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_830 = _T_11 ? _GEN_302 : REG__6_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_831 = _T_11 ? _GEN_303 : REG__7_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_832 = _T_11 ? _GEN_304 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_833 = _T_11 ? _GEN_305 : REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_834 = _T_11 ? _GEN_306 : REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_835 = _T_11 ? _GEN_307 : REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_836 = _T_11 ? _GEN_308 : REG__4_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_837 = _T_11 ? _GEN_309 : REG__5_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_838 = _T_11 ? _GEN_310 : REG__6_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_839 = _T_11 ? _GEN_311 : REG__7_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_840 = _T_11 ? _GEN_312 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_841 = _T_11 ? _GEN_313 : REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_842 = _T_11 ? _GEN_314 : REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_843 = _T_11 ? _GEN_315 : REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_844 = _T_11 ? _GEN_316 : REG__4_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_845 = _T_11 ? _GEN_317 : REG__5_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_846 = _T_11 ? _GEN_318 : REG__6_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_847 = _T_11 ? _GEN_319 : REG__7_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_848 = _T_11 ? _GEN_320 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_849 = _T_11 ? _GEN_321 : REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_850 = _T_11 ? _GEN_322 : REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_851 = _T_11 ? _GEN_323 : REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_852 = _T_11 ? _GEN_324 : REG__4_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_853 = _T_11 ? _GEN_325 : REG__5_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_854 = _T_11 ? _GEN_326 : REG__6_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_855 = _T_11 ? _GEN_327 : REG__7_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_856 = _T_11 ? _GEN_328 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_857 = _T_11 ? _GEN_329 : REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_858 = _T_11 ? _GEN_330 : REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_859 = _T_11 ? _GEN_331 : REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_860 = _T_11 ? _GEN_332 : REG__4_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_861 = _T_11 ? _GEN_333 : REG__5_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_862 = _T_11 ? _GEN_334 : REG__6_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_863 = _T_11 ? _GEN_335 : REG__7_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_864 = _T_11 ? _GEN_336 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_865 = _T_11 ? _GEN_337 : REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_866 = _T_11 ? _GEN_338 : REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_867 = _T_11 ? _GEN_339 : REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_868 = _T_11 ? _GEN_340 : REG__4_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_869 = _T_11 ? _GEN_341 : REG__5_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_870 = _T_11 ? _GEN_342 : REG__6_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_871 = _T_11 ? _GEN_343 : REG__7_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_872 = _T_11 ? _GEN_344 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_873 = _T_11 ? _GEN_345 : REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_874 = _T_11 ? _GEN_346 : REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_875 = _T_11 ? _GEN_347 : REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_876 = _T_11 ? _GEN_348 : REG__4_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_877 = _T_11 ? _GEN_349 : REG__5_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_878 = _T_11 ? _GEN_350 : REG__6_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_879 = _T_11 ? _GEN_351 : REG__7_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_888 = _T_11 ? _GEN_360 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_889 = _T_11 ? _GEN_361 : REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_890 = _T_11 ? _GEN_362 : REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_891 = _T_11 ? _GEN_363 : REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_892 = _T_11 ? _GEN_364 : REG__4_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_893 = _T_11 ? _GEN_365 : REG__5_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_894 = _T_11 ? _GEN_366 : REG__6_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_895 = _T_11 ? _GEN_367 : REG__7_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_896 = _T_11 ? _GEN_368 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_897 = _T_11 ? _GEN_369 : REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_898 = _T_11 ? _GEN_370 : REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_899 = _T_11 ? _GEN_371 : REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_900 = _T_11 ? _GEN_372 : REG__4_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_901 = _T_11 ? _GEN_373 : REG__5_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_902 = _T_11 ? _GEN_374 : REG__6_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_903 = _T_11 ? _GEN_375 : REG__7_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_976 = _T_11 ? _GEN_448 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_977 = _T_11 ? _GEN_449 : REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_978 = _T_11 ? _GEN_450 : REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_979 = _T_11 ? _GEN_451 : REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_980 = _T_11 ? _GEN_452 : REG__4_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_981 = _T_11 ? _GEN_453 : REG__5_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_982 = _T_11 ? _GEN_454 : REG__6_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_983 = _T_11 ? _GEN_455 : REG__7_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1032 = _T_11 ? _GEN_504 : REG__0_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1033 = _T_11 ? _GEN_505 : REG__1_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1034 = _T_11 ? _GEN_506 : REG__2_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1035 = _T_11 ? _GEN_507 : REG__3_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1036 = _T_11 ? _GEN_508 : REG__4_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1037 = _T_11 ? _GEN_509 : REG__5_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1038 = _T_11 ? _GEN_510 : REG__6_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1039 = _T_11 ? _GEN_511 : REG__7_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1040 = _T_11 ? _GEN_512 : REG__0_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1041 = _T_11 ? _GEN_513 : REG__1_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1042 = _T_11 ? _GEN_514 : REG__2_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1043 = _T_11 ? _GEN_515 : REG__3_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1044 = _T_11 ? _GEN_516 : REG__4_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1045 = _T_11 ? _GEN_517 : REG__5_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1046 = _T_11 ? _GEN_518 : REG__6_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1047 = _T_11 ? _GEN_519 : REG__7_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1048 = _T_11 ? _GEN_520 : REG__0_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1049 = _T_11 ? _GEN_521 : REG__1_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1050 = _T_11 ? _GEN_522 : REG__2_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1051 = _T_11 ? _GEN_523 : REG__3_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1052 = _T_11 ? _GEN_524 : REG__4_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1053 = _T_11 ? _GEN_525 : REG__5_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1054 = _T_11 ? _GEN_526 : REG__6_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1055 = _T_11 ? _GEN_527 : REG__7_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _T_20 = 3'h1 + REG_1; // @[PipelineVector.scala 46:45]
  wire [2:0] _GEN_3716 = {{1'd0}, _T_10}; // @[PipelineVector.scala 47:42]
  wire [2:0] _T_22 = REG_1 + _GEN_3716; // @[PipelineVector.scala 47:42]
  wire [63:0] _GEN_2666 = 3'h1 == REG_2 ? REG__1_data_imm : REG__0_data_imm; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2667 = 3'h2 == REG_2 ? REG__2_data_imm : _GEN_2666; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2668 = 3'h3 == REG_2 ? REG__3_data_imm : _GEN_2667; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2669 = 3'h4 == REG_2 ? REG__4_data_imm : _GEN_2668; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2670 = 3'h5 == REG_2 ? REG__5_data_imm : _GEN_2669; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2671 = 3'h6 == REG_2 ? REG__6_data_imm : _GEN_2670; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2698 = 3'h1 == REG_2 ? REG__1_ctrl_isMou : REG__0_ctrl_isMou; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2699 = 3'h2 == REG_2 ? REG__2_ctrl_isMou : _GEN_2698; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2700 = 3'h3 == REG_2 ? REG__3_ctrl_isMou : _GEN_2699; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2701 = 3'h4 == REG_2 ? REG__4_ctrl_isMou : _GEN_2700; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2702 = 3'h5 == REG_2 ? REG__5_ctrl_isMou : _GEN_2701; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2703 = 3'h6 == REG_2 ? REG__6_ctrl_isMou : _GEN_2702; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2754 = 3'h1 == REG_2 ? REG__1_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2755 = 3'h2 == REG_2 ? REG__2_ctrl_rfDest : _GEN_2754; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2756 = 3'h3 == REG_2 ? REG__3_ctrl_rfDest : _GEN_2755; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2757 = 3'h4 == REG_2 ? REG__4_ctrl_rfDest : _GEN_2756; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2758 = 3'h5 == REG_2 ? REG__5_ctrl_rfDest : _GEN_2757; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2759 = 3'h6 == REG_2 ? REG__6_ctrl_rfDest : _GEN_2758; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2762 = 3'h1 == REG_2 ? REG__1_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2763 = 3'h2 == REG_2 ? REG__2_ctrl_rfWen : _GEN_2762; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2764 = 3'h3 == REG_2 ? REG__3_ctrl_rfWen : _GEN_2763; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2765 = 3'h4 == REG_2 ? REG__4_ctrl_rfWen : _GEN_2764; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2766 = 3'h5 == REG_2 ? REG__5_ctrl_rfWen : _GEN_2765; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2767 = 3'h6 == REG_2 ? REG__6_ctrl_rfWen : _GEN_2766; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2770 = 3'h1 == REG_2 ? REG__1_ctrl_rfSrc3 : REG__0_ctrl_rfSrc3; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2771 = 3'h2 == REG_2 ? REG__2_ctrl_rfSrc3 : _GEN_2770; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2772 = 3'h3 == REG_2 ? REG__3_ctrl_rfSrc3 : _GEN_2771; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2773 = 3'h4 == REG_2 ? REG__4_ctrl_rfSrc3 : _GEN_2772; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2774 = 3'h5 == REG_2 ? REG__5_ctrl_rfSrc3 : _GEN_2773; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2775 = 3'h6 == REG_2 ? REG__6_ctrl_rfSrc3 : _GEN_2774; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2778 = 3'h1 == REG_2 ? REG__1_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2779 = 3'h2 == REG_2 ? REG__2_ctrl_rfSrc2 : _GEN_2778; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2780 = 3'h3 == REG_2 ? REG__3_ctrl_rfSrc2 : _GEN_2779; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2781 = 3'h4 == REG_2 ? REG__4_ctrl_rfSrc2 : _GEN_2780; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2782 = 3'h5 == REG_2 ? REG__5_ctrl_rfSrc2 : _GEN_2781; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2783 = 3'h6 == REG_2 ? REG__6_ctrl_rfSrc2 : _GEN_2782; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2786 = 3'h1 == REG_2 ? REG__1_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2787 = 3'h2 == REG_2 ? REG__2_ctrl_rfSrc1 : _GEN_2786; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2788 = 3'h3 == REG_2 ? REG__3_ctrl_rfSrc1 : _GEN_2787; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2789 = 3'h4 == REG_2 ? REG__4_ctrl_rfSrc1 : _GEN_2788; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2790 = 3'h5 == REG_2 ? REG__5_ctrl_rfSrc1 : _GEN_2789; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2791 = 3'h6 == REG_2 ? REG__6_ctrl_rfSrc1 : _GEN_2790; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2794 = 3'h1 == REG_2 ? REG__1_ctrl_func23 : REG__0_ctrl_func23; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2795 = 3'h2 == REG_2 ? REG__2_ctrl_func23 : _GEN_2794; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2796 = 3'h3 == REG_2 ? REG__3_ctrl_func23 : _GEN_2795; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2797 = 3'h4 == REG_2 ? REG__4_ctrl_func23 : _GEN_2796; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2798 = 3'h5 == REG_2 ? REG__5_ctrl_func23 : _GEN_2797; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2799 = 3'h6 == REG_2 ? REG__6_ctrl_func23 : _GEN_2798; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2802 = 3'h1 == REG_2 ? REG__1_ctrl_func24 : REG__0_ctrl_func24; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2803 = 3'h2 == REG_2 ? REG__2_ctrl_func24 : _GEN_2802; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2804 = 3'h3 == REG_2 ? REG__3_ctrl_func24 : _GEN_2803; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2805 = 3'h4 == REG_2 ? REG__4_ctrl_func24 : _GEN_2804; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2806 = 3'h5 == REG_2 ? REG__5_ctrl_func24 : _GEN_2805; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2807 = 3'h6 == REG_2 ? REG__6_ctrl_func24 : _GEN_2806; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_2810 = 3'h1 == REG_2 ? REG__1_ctrl_funct3 : REG__0_ctrl_funct3; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_2811 = 3'h2 == REG_2 ? REG__2_ctrl_funct3 : _GEN_2810; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_2812 = 3'h3 == REG_2 ? REG__3_ctrl_funct3 : _GEN_2811; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_2813 = 3'h4 == REG_2 ? REG__4_ctrl_funct3 : _GEN_2812; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_2814 = 3'h5 == REG_2 ? REG__5_ctrl_funct3 : _GEN_2813; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_2815 = 3'h6 == REG_2 ? REG__6_ctrl_funct3 : _GEN_2814; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_2818 = 3'h1 == REG_2 ? REG__1_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_2819 = 3'h2 == REG_2 ? REG__2_ctrl_fuOpType : _GEN_2818; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_2820 = 3'h3 == REG_2 ? REG__3_ctrl_fuOpType : _GEN_2819; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_2821 = 3'h4 == REG_2 ? REG__4_ctrl_fuOpType : _GEN_2820; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_2822 = 3'h5 == REG_2 ? REG__5_ctrl_fuOpType : _GEN_2821; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_2823 = 3'h6 == REG_2 ? REG__6_ctrl_fuOpType : _GEN_2822; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2826 = 3'h1 == REG_2 ? REG__1_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2827 = 3'h2 == REG_2 ? REG__2_ctrl_fuType : _GEN_2826; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2828 = 3'h3 == REG_2 ? REG__3_ctrl_fuType : _GEN_2827; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2829 = 3'h4 == REG_2 ? REG__4_ctrl_fuType : _GEN_2828; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2830 = 3'h5 == REG_2 ? REG__5_ctrl_fuType : _GEN_2829; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2831 = 3'h6 == REG_2 ? REG__6_ctrl_fuType : _GEN_2830; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2834 = 3'h1 == REG_2 ? REG__1_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2835 = 3'h2 == REG_2 ? REG__2_ctrl_src2Type : _GEN_2834; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2836 = 3'h3 == REG_2 ? REG__3_ctrl_src2Type : _GEN_2835; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2837 = 3'h4 == REG_2 ? REG__4_ctrl_src2Type : _GEN_2836; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2838 = 3'h5 == REG_2 ? REG__5_ctrl_src2Type : _GEN_2837; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2839 = 3'h6 == REG_2 ? REG__6_ctrl_src2Type : _GEN_2838; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2842 = 3'h1 == REG_2 ? REG__1_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2843 = 3'h2 == REG_2 ? REG__2_ctrl_src1Type : _GEN_2842; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2844 = 3'h3 == REG_2 ? REG__3_ctrl_src1Type : _GEN_2843; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2845 = 3'h4 == REG_2 ? REG__4_ctrl_src1Type : _GEN_2844; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2846 = 3'h5 == REG_2 ? REG__5_ctrl_src1Type : _GEN_2845; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2847 = 3'h6 == REG_2 ? REG__6_ctrl_src1Type : _GEN_2846; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2850 = 3'h1 == REG_2 ? REG__1_cf_instrType : REG__0_cf_instrType; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2851 = 3'h2 == REG_2 ? REG__2_cf_instrType : _GEN_2850; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2852 = 3'h3 == REG_2 ? REG__3_cf_instrType : _GEN_2851; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2853 = 3'h4 == REG_2 ? REG__4_cf_instrType : _GEN_2852; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2854 = 3'h5 == REG_2 ? REG__5_cf_instrType : _GEN_2853; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_2855 = 3'h6 == REG_2 ? REG__6_cf_instrType : _GEN_2854; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2866 = 3'h1 == REG_2 ? REG__1_cf_runahead_checkpoint_id : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2867 = 3'h2 == REG_2 ? REG__2_cf_runahead_checkpoint_id : _GEN_2866; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2868 = 3'h3 == REG_2 ? REG__3_cf_runahead_checkpoint_id : _GEN_2867; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2869 = 3'h4 == REG_2 ? REG__4_cf_runahead_checkpoint_id : _GEN_2868; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2870 = 3'h5 == REG_2 ? REG__5_cf_runahead_checkpoint_id : _GEN_2869; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_2871 = 3'h6 == REG_2 ? REG__6_cf_runahead_checkpoint_id : _GEN_2870; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2874 = 3'h1 == REG_2 ? REG__1_cf_crossPageIPFFix : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2875 = 3'h2 == REG_2 ? REG__2_cf_crossPageIPFFix : _GEN_2874; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2876 = 3'h3 == REG_2 ? REG__3_cf_crossPageIPFFix : _GEN_2875; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2877 = 3'h4 == REG_2 ? REG__4_cf_crossPageIPFFix : _GEN_2876; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2878 = 3'h5 == REG_2 ? REG__5_cf_crossPageIPFFix : _GEN_2877; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2879 = 3'h6 == REG_2 ? REG__6_cf_crossPageIPFFix : _GEN_2878; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2890 = 3'h1 == REG_2 ? REG__1_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2891 = 3'h2 == REG_2 ? REG__2_cf_brIdx : _GEN_2890; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2892 = 3'h3 == REG_2 ? REG__3_cf_brIdx : _GEN_2891; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2893 = 3'h4 == REG_2 ? REG__4_cf_brIdx : _GEN_2892; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2894 = 3'h5 == REG_2 ? REG__5_cf_brIdx : _GEN_2893; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_2895 = 3'h6 == REG_2 ? REG__6_cf_brIdx : _GEN_2894; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2898 = 3'h1 == REG_2 ? REG__1_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2899 = 3'h2 == REG_2 ? REG__2_cf_intrVec_0 : _GEN_2898; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2900 = 3'h3 == REG_2 ? REG__3_cf_intrVec_0 : _GEN_2899; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2901 = 3'h4 == REG_2 ? REG__4_cf_intrVec_0 : _GEN_2900; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2902 = 3'h5 == REG_2 ? REG__5_cf_intrVec_0 : _GEN_2901; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2903 = 3'h6 == REG_2 ? REG__6_cf_intrVec_0 : _GEN_2902; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2906 = 3'h1 == REG_2 ? REG__1_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2907 = 3'h2 == REG_2 ? REG__2_cf_intrVec_1 : _GEN_2906; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2908 = 3'h3 == REG_2 ? REG__3_cf_intrVec_1 : _GEN_2907; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2909 = 3'h4 == REG_2 ? REG__4_cf_intrVec_1 : _GEN_2908; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2910 = 3'h5 == REG_2 ? REG__5_cf_intrVec_1 : _GEN_2909; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2911 = 3'h6 == REG_2 ? REG__6_cf_intrVec_1 : _GEN_2910; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2914 = 3'h1 == REG_2 ? REG__1_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2915 = 3'h2 == REG_2 ? REG__2_cf_intrVec_2 : _GEN_2914; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2916 = 3'h3 == REG_2 ? REG__3_cf_intrVec_2 : _GEN_2915; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2917 = 3'h4 == REG_2 ? REG__4_cf_intrVec_2 : _GEN_2916; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2918 = 3'h5 == REG_2 ? REG__5_cf_intrVec_2 : _GEN_2917; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2919 = 3'h6 == REG_2 ? REG__6_cf_intrVec_2 : _GEN_2918; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2922 = 3'h1 == REG_2 ? REG__1_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2923 = 3'h2 == REG_2 ? REG__2_cf_intrVec_3 : _GEN_2922; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2924 = 3'h3 == REG_2 ? REG__3_cf_intrVec_3 : _GEN_2923; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2925 = 3'h4 == REG_2 ? REG__4_cf_intrVec_3 : _GEN_2924; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2926 = 3'h5 == REG_2 ? REG__5_cf_intrVec_3 : _GEN_2925; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2927 = 3'h6 == REG_2 ? REG__6_cf_intrVec_3 : _GEN_2926; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2930 = 3'h1 == REG_2 ? REG__1_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2931 = 3'h2 == REG_2 ? REG__2_cf_intrVec_4 : _GEN_2930; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2932 = 3'h3 == REG_2 ? REG__3_cf_intrVec_4 : _GEN_2931; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2933 = 3'h4 == REG_2 ? REG__4_cf_intrVec_4 : _GEN_2932; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2934 = 3'h5 == REG_2 ? REG__5_cf_intrVec_4 : _GEN_2933; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2935 = 3'h6 == REG_2 ? REG__6_cf_intrVec_4 : _GEN_2934; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2938 = 3'h1 == REG_2 ? REG__1_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2939 = 3'h2 == REG_2 ? REG__2_cf_intrVec_5 : _GEN_2938; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2940 = 3'h3 == REG_2 ? REG__3_cf_intrVec_5 : _GEN_2939; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2941 = 3'h4 == REG_2 ? REG__4_cf_intrVec_5 : _GEN_2940; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2942 = 3'h5 == REG_2 ? REG__5_cf_intrVec_5 : _GEN_2941; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2943 = 3'h6 == REG_2 ? REG__6_cf_intrVec_5 : _GEN_2942; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2946 = 3'h1 == REG_2 ? REG__1_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2947 = 3'h2 == REG_2 ? REG__2_cf_intrVec_6 : _GEN_2946; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2948 = 3'h3 == REG_2 ? REG__3_cf_intrVec_6 : _GEN_2947; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2949 = 3'h4 == REG_2 ? REG__4_cf_intrVec_6 : _GEN_2948; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2950 = 3'h5 == REG_2 ? REG__5_cf_intrVec_6 : _GEN_2949; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2951 = 3'h6 == REG_2 ? REG__6_cf_intrVec_6 : _GEN_2950; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2954 = 3'h1 == REG_2 ? REG__1_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2955 = 3'h2 == REG_2 ? REG__2_cf_intrVec_7 : _GEN_2954; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2956 = 3'h3 == REG_2 ? REG__3_cf_intrVec_7 : _GEN_2955; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2957 = 3'h4 == REG_2 ? REG__4_cf_intrVec_7 : _GEN_2956; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2958 = 3'h5 == REG_2 ? REG__5_cf_intrVec_7 : _GEN_2957; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2959 = 3'h6 == REG_2 ? REG__6_cf_intrVec_7 : _GEN_2958; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2962 = 3'h1 == REG_2 ? REG__1_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2963 = 3'h2 == REG_2 ? REG__2_cf_intrVec_8 : _GEN_2962; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2964 = 3'h3 == REG_2 ? REG__3_cf_intrVec_8 : _GEN_2963; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2965 = 3'h4 == REG_2 ? REG__4_cf_intrVec_8 : _GEN_2964; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2966 = 3'h5 == REG_2 ? REG__5_cf_intrVec_8 : _GEN_2965; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2967 = 3'h6 == REG_2 ? REG__6_cf_intrVec_8 : _GEN_2966; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2970 = 3'h1 == REG_2 ? REG__1_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2971 = 3'h2 == REG_2 ? REG__2_cf_intrVec_9 : _GEN_2970; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2972 = 3'h3 == REG_2 ? REG__3_cf_intrVec_9 : _GEN_2971; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2973 = 3'h4 == REG_2 ? REG__4_cf_intrVec_9 : _GEN_2972; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2974 = 3'h5 == REG_2 ? REG__5_cf_intrVec_9 : _GEN_2973; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2975 = 3'h6 == REG_2 ? REG__6_cf_intrVec_9 : _GEN_2974; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2978 = 3'h1 == REG_2 ? REG__1_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2979 = 3'h2 == REG_2 ? REG__2_cf_intrVec_10 : _GEN_2978; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2980 = 3'h3 == REG_2 ? REG__3_cf_intrVec_10 : _GEN_2979; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2981 = 3'h4 == REG_2 ? REG__4_cf_intrVec_10 : _GEN_2980; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2982 = 3'h5 == REG_2 ? REG__5_cf_intrVec_10 : _GEN_2981; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2983 = 3'h6 == REG_2 ? REG__6_cf_intrVec_10 : _GEN_2982; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2986 = 3'h1 == REG_2 ? REG__1_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2987 = 3'h2 == REG_2 ? REG__2_cf_intrVec_11 : _GEN_2986; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2988 = 3'h3 == REG_2 ? REG__3_cf_intrVec_11 : _GEN_2987; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2989 = 3'h4 == REG_2 ? REG__4_cf_intrVec_11 : _GEN_2988; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2990 = 3'h5 == REG_2 ? REG__5_cf_intrVec_11 : _GEN_2989; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_2991 = 3'h6 == REG_2 ? REG__6_cf_intrVec_11 : _GEN_2990; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3002 = 3'h1 == REG_2 ? REG__1_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3003 = 3'h2 == REG_2 ? REG__2_cf_exceptionVec_1 : _GEN_3002; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3004 = 3'h3 == REG_2 ? REG__3_cf_exceptionVec_1 : _GEN_3003; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3005 = 3'h4 == REG_2 ? REG__4_cf_exceptionVec_1 : _GEN_3004; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3006 = 3'h5 == REG_2 ? REG__5_cf_exceptionVec_1 : _GEN_3005; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3007 = 3'h6 == REG_2 ? REG__6_cf_exceptionVec_1 : _GEN_3006; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3010 = 3'h1 == REG_2 ? REG__1_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3011 = 3'h2 == REG_2 ? REG__2_cf_exceptionVec_2 : _GEN_3010; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3012 = 3'h3 == REG_2 ? REG__3_cf_exceptionVec_2 : _GEN_3011; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3013 = 3'h4 == REG_2 ? REG__4_cf_exceptionVec_2 : _GEN_3012; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3014 = 3'h5 == REG_2 ? REG__5_cf_exceptionVec_2 : _GEN_3013; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3015 = 3'h6 == REG_2 ? REG__6_cf_exceptionVec_2 : _GEN_3014; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3090 = 3'h1 == REG_2 ? REG__1_cf_exceptionVec_12 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3091 = 3'h2 == REG_2 ? REG__2_cf_exceptionVec_12 : _GEN_3090; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3092 = 3'h3 == REG_2 ? REG__3_cf_exceptionVec_12 : _GEN_3091; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3093 = 3'h4 == REG_2 ? REG__4_cf_exceptionVec_12 : _GEN_3092; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3094 = 3'h5 == REG_2 ? REG__5_cf_exceptionVec_12 : _GEN_3093; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_3095 = 3'h6 == REG_2 ? REG__6_cf_exceptionVec_12 : _GEN_3094; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3146 = 3'h1 == REG_2 ? REG__1_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3147 = 3'h2 == REG_2 ? REG__2_cf_pnpc : _GEN_3146; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3148 = 3'h3 == REG_2 ? REG__3_cf_pnpc : _GEN_3147; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3149 = 3'h4 == REG_2 ? REG__4_cf_pnpc : _GEN_3148; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3150 = 3'h5 == REG_2 ? REG__5_cf_pnpc : _GEN_3149; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3151 = 3'h6 == REG_2 ? REG__6_cf_pnpc : _GEN_3150; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3154 = 3'h1 == REG_2 ? REG__1_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3155 = 3'h2 == REG_2 ? REG__2_cf_pc : _GEN_3154; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3156 = 3'h3 == REG_2 ? REG__3_cf_pc : _GEN_3155; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3157 = 3'h4 == REG_2 ? REG__4_cf_pc : _GEN_3156; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3158 = 3'h5 == REG_2 ? REG__5_cf_pc : _GEN_3157; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_3159 = 3'h6 == REG_2 ? REG__6_cf_pc : _GEN_3158; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_3162 = 3'h1 == REG_2 ? REG__1_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_3163 = 3'h2 == REG_2 ? REG__2_cf_instr : _GEN_3162; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_3164 = 3'h3 == REG_2 ? REG__3_cf_instr : _GEN_3163; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_3165 = 3'h4 == REG_2 ? REG__4_cf_instr : _GEN_3164; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_3166 = 3'h5 == REG_2 ? REG__5_cf_instr : _GEN_3165; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_3167 = 3'h6 == REG_2 ? REG__6_cf_instr : _GEN_3166; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _T_29 = REG_2 + 3'h1; // @[PipelineVector.scala 59:42]
  wire [63:0] _GEN_3194 = 3'h1 == _T_29 ? REG__1_data_imm : REG__0_data_imm; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3195 = 3'h2 == _T_29 ? REG__2_data_imm : _GEN_3194; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3196 = 3'h3 == _T_29 ? REG__3_data_imm : _GEN_3195; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3197 = 3'h4 == _T_29 ? REG__4_data_imm : _GEN_3196; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3198 = 3'h5 == _T_29 ? REG__5_data_imm : _GEN_3197; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3199 = 3'h6 == _T_29 ? REG__6_data_imm : _GEN_3198; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3226 = 3'h1 == _T_29 ? REG__1_ctrl_isMou : REG__0_ctrl_isMou; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3227 = 3'h2 == _T_29 ? REG__2_ctrl_isMou : _GEN_3226; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3228 = 3'h3 == _T_29 ? REG__3_ctrl_isMou : _GEN_3227; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3229 = 3'h4 == _T_29 ? REG__4_ctrl_isMou : _GEN_3228; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3230 = 3'h5 == _T_29 ? REG__5_ctrl_isMou : _GEN_3229; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3231 = 3'h6 == _T_29 ? REG__6_ctrl_isMou : _GEN_3230; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3282 = 3'h1 == _T_29 ? REG__1_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3283 = 3'h2 == _T_29 ? REG__2_ctrl_rfDest : _GEN_3282; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3284 = 3'h3 == _T_29 ? REG__3_ctrl_rfDest : _GEN_3283; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3285 = 3'h4 == _T_29 ? REG__4_ctrl_rfDest : _GEN_3284; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3286 = 3'h5 == _T_29 ? REG__5_ctrl_rfDest : _GEN_3285; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3287 = 3'h6 == _T_29 ? REG__6_ctrl_rfDest : _GEN_3286; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3290 = 3'h1 == _T_29 ? REG__1_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3291 = 3'h2 == _T_29 ? REG__2_ctrl_rfWen : _GEN_3290; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3292 = 3'h3 == _T_29 ? REG__3_ctrl_rfWen : _GEN_3291; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3293 = 3'h4 == _T_29 ? REG__4_ctrl_rfWen : _GEN_3292; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3294 = 3'h5 == _T_29 ? REG__5_ctrl_rfWen : _GEN_3293; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3295 = 3'h6 == _T_29 ? REG__6_ctrl_rfWen : _GEN_3294; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3298 = 3'h1 == _T_29 ? REG__1_ctrl_rfSrc3 : REG__0_ctrl_rfSrc3; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3299 = 3'h2 == _T_29 ? REG__2_ctrl_rfSrc3 : _GEN_3298; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3300 = 3'h3 == _T_29 ? REG__3_ctrl_rfSrc3 : _GEN_3299; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3301 = 3'h4 == _T_29 ? REG__4_ctrl_rfSrc3 : _GEN_3300; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3302 = 3'h5 == _T_29 ? REG__5_ctrl_rfSrc3 : _GEN_3301; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3303 = 3'h6 == _T_29 ? REG__6_ctrl_rfSrc3 : _GEN_3302; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3306 = 3'h1 == _T_29 ? REG__1_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3307 = 3'h2 == _T_29 ? REG__2_ctrl_rfSrc2 : _GEN_3306; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3308 = 3'h3 == _T_29 ? REG__3_ctrl_rfSrc2 : _GEN_3307; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3309 = 3'h4 == _T_29 ? REG__4_ctrl_rfSrc2 : _GEN_3308; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3310 = 3'h5 == _T_29 ? REG__5_ctrl_rfSrc2 : _GEN_3309; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3311 = 3'h6 == _T_29 ? REG__6_ctrl_rfSrc2 : _GEN_3310; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3314 = 3'h1 == _T_29 ? REG__1_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3315 = 3'h2 == _T_29 ? REG__2_ctrl_rfSrc1 : _GEN_3314; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3316 = 3'h3 == _T_29 ? REG__3_ctrl_rfSrc1 : _GEN_3315; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3317 = 3'h4 == _T_29 ? REG__4_ctrl_rfSrc1 : _GEN_3316; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3318 = 3'h5 == _T_29 ? REG__5_ctrl_rfSrc1 : _GEN_3317; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3319 = 3'h6 == _T_29 ? REG__6_ctrl_rfSrc1 : _GEN_3318; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3322 = 3'h1 == _T_29 ? REG__1_ctrl_func23 : REG__0_ctrl_func23; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3323 = 3'h2 == _T_29 ? REG__2_ctrl_func23 : _GEN_3322; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3324 = 3'h3 == _T_29 ? REG__3_ctrl_func23 : _GEN_3323; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3325 = 3'h4 == _T_29 ? REG__4_ctrl_func23 : _GEN_3324; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3326 = 3'h5 == _T_29 ? REG__5_ctrl_func23 : _GEN_3325; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3327 = 3'h6 == _T_29 ? REG__6_ctrl_func23 : _GEN_3326; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3330 = 3'h1 == _T_29 ? REG__1_ctrl_func24 : REG__0_ctrl_func24; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3331 = 3'h2 == _T_29 ? REG__2_ctrl_func24 : _GEN_3330; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3332 = 3'h3 == _T_29 ? REG__3_ctrl_func24 : _GEN_3331; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3333 = 3'h4 == _T_29 ? REG__4_ctrl_func24 : _GEN_3332; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3334 = 3'h5 == _T_29 ? REG__5_ctrl_func24 : _GEN_3333; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3335 = 3'h6 == _T_29 ? REG__6_ctrl_func24 : _GEN_3334; // @[PipelineVector.scala 60:{15,15}]
  wire [2:0] _GEN_3338 = 3'h1 == _T_29 ? REG__1_ctrl_funct3 : REG__0_ctrl_funct3; // @[PipelineVector.scala 60:{15,15}]
  wire [2:0] _GEN_3339 = 3'h2 == _T_29 ? REG__2_ctrl_funct3 : _GEN_3338; // @[PipelineVector.scala 60:{15,15}]
  wire [2:0] _GEN_3340 = 3'h3 == _T_29 ? REG__3_ctrl_funct3 : _GEN_3339; // @[PipelineVector.scala 60:{15,15}]
  wire [2:0] _GEN_3341 = 3'h4 == _T_29 ? REG__4_ctrl_funct3 : _GEN_3340; // @[PipelineVector.scala 60:{15,15}]
  wire [2:0] _GEN_3342 = 3'h5 == _T_29 ? REG__5_ctrl_funct3 : _GEN_3341; // @[PipelineVector.scala 60:{15,15}]
  wire [2:0] _GEN_3343 = 3'h6 == _T_29 ? REG__6_ctrl_funct3 : _GEN_3342; // @[PipelineVector.scala 60:{15,15}]
  wire [6:0] _GEN_3346 = 3'h1 == _T_29 ? REG__1_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 60:{15,15}]
  wire [6:0] _GEN_3347 = 3'h2 == _T_29 ? REG__2_ctrl_fuOpType : _GEN_3346; // @[PipelineVector.scala 60:{15,15}]
  wire [6:0] _GEN_3348 = 3'h3 == _T_29 ? REG__3_ctrl_fuOpType : _GEN_3347; // @[PipelineVector.scala 60:{15,15}]
  wire [6:0] _GEN_3349 = 3'h4 == _T_29 ? REG__4_ctrl_fuOpType : _GEN_3348; // @[PipelineVector.scala 60:{15,15}]
  wire [6:0] _GEN_3350 = 3'h5 == _T_29 ? REG__5_ctrl_fuOpType : _GEN_3349; // @[PipelineVector.scala 60:{15,15}]
  wire [6:0] _GEN_3351 = 3'h6 == _T_29 ? REG__6_ctrl_fuOpType : _GEN_3350; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3354 = 3'h1 == _T_29 ? REG__1_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3355 = 3'h2 == _T_29 ? REG__2_ctrl_fuType : _GEN_3354; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3356 = 3'h3 == _T_29 ? REG__3_ctrl_fuType : _GEN_3355; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3357 = 3'h4 == _T_29 ? REG__4_ctrl_fuType : _GEN_3356; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3358 = 3'h5 == _T_29 ? REG__5_ctrl_fuType : _GEN_3357; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3359 = 3'h6 == _T_29 ? REG__6_ctrl_fuType : _GEN_3358; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3362 = 3'h1 == _T_29 ? REG__1_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3363 = 3'h2 == _T_29 ? REG__2_ctrl_src2Type : _GEN_3362; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3364 = 3'h3 == _T_29 ? REG__3_ctrl_src2Type : _GEN_3363; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3365 = 3'h4 == _T_29 ? REG__4_ctrl_src2Type : _GEN_3364; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3366 = 3'h5 == _T_29 ? REG__5_ctrl_src2Type : _GEN_3365; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3367 = 3'h6 == _T_29 ? REG__6_ctrl_src2Type : _GEN_3366; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3370 = 3'h1 == _T_29 ? REG__1_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3371 = 3'h2 == _T_29 ? REG__2_ctrl_src1Type : _GEN_3370; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3372 = 3'h3 == _T_29 ? REG__3_ctrl_src1Type : _GEN_3371; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3373 = 3'h4 == _T_29 ? REG__4_ctrl_src1Type : _GEN_3372; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3374 = 3'h5 == _T_29 ? REG__5_ctrl_src1Type : _GEN_3373; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3375 = 3'h6 == _T_29 ? REG__6_ctrl_src1Type : _GEN_3374; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3378 = 3'h1 == _T_29 ? REG__1_cf_instrType : REG__0_cf_instrType; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3379 = 3'h2 == _T_29 ? REG__2_cf_instrType : _GEN_3378; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3380 = 3'h3 == _T_29 ? REG__3_cf_instrType : _GEN_3379; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3381 = 3'h4 == _T_29 ? REG__4_cf_instrType : _GEN_3380; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3382 = 3'h5 == _T_29 ? REG__5_cf_instrType : _GEN_3381; // @[PipelineVector.scala 60:{15,15}]
  wire [4:0] _GEN_3383 = 3'h6 == _T_29 ? REG__6_cf_instrType : _GEN_3382; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3394 = 3'h1 == _T_29 ? REG__1_cf_runahead_checkpoint_id : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3395 = 3'h2 == _T_29 ? REG__2_cf_runahead_checkpoint_id : _GEN_3394; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3396 = 3'h3 == _T_29 ? REG__3_cf_runahead_checkpoint_id : _GEN_3395; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3397 = 3'h4 == _T_29 ? REG__4_cf_runahead_checkpoint_id : _GEN_3396; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3398 = 3'h5 == _T_29 ? REG__5_cf_runahead_checkpoint_id : _GEN_3397; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3399 = 3'h6 == _T_29 ? REG__6_cf_runahead_checkpoint_id : _GEN_3398; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3402 = 3'h1 == _T_29 ? REG__1_cf_crossPageIPFFix : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3403 = 3'h2 == _T_29 ? REG__2_cf_crossPageIPFFix : _GEN_3402; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3404 = 3'h3 == _T_29 ? REG__3_cf_crossPageIPFFix : _GEN_3403; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3405 = 3'h4 == _T_29 ? REG__4_cf_crossPageIPFFix : _GEN_3404; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3406 = 3'h5 == _T_29 ? REG__5_cf_crossPageIPFFix : _GEN_3405; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3407 = 3'h6 == _T_29 ? REG__6_cf_crossPageIPFFix : _GEN_3406; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3418 = 3'h1 == _T_29 ? REG__1_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3419 = 3'h2 == _T_29 ? REG__2_cf_brIdx : _GEN_3418; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3420 = 3'h3 == _T_29 ? REG__3_cf_brIdx : _GEN_3419; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3421 = 3'h4 == _T_29 ? REG__4_cf_brIdx : _GEN_3420; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3422 = 3'h5 == _T_29 ? REG__5_cf_brIdx : _GEN_3421; // @[PipelineVector.scala 60:{15,15}]
  wire [3:0] _GEN_3423 = 3'h6 == _T_29 ? REG__6_cf_brIdx : _GEN_3422; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3426 = 3'h1 == _T_29 ? REG__1_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3427 = 3'h2 == _T_29 ? REG__2_cf_intrVec_0 : _GEN_3426; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3428 = 3'h3 == _T_29 ? REG__3_cf_intrVec_0 : _GEN_3427; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3429 = 3'h4 == _T_29 ? REG__4_cf_intrVec_0 : _GEN_3428; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3430 = 3'h5 == _T_29 ? REG__5_cf_intrVec_0 : _GEN_3429; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3431 = 3'h6 == _T_29 ? REG__6_cf_intrVec_0 : _GEN_3430; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3434 = 3'h1 == _T_29 ? REG__1_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3435 = 3'h2 == _T_29 ? REG__2_cf_intrVec_1 : _GEN_3434; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3436 = 3'h3 == _T_29 ? REG__3_cf_intrVec_1 : _GEN_3435; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3437 = 3'h4 == _T_29 ? REG__4_cf_intrVec_1 : _GEN_3436; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3438 = 3'h5 == _T_29 ? REG__5_cf_intrVec_1 : _GEN_3437; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3439 = 3'h6 == _T_29 ? REG__6_cf_intrVec_1 : _GEN_3438; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3442 = 3'h1 == _T_29 ? REG__1_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3443 = 3'h2 == _T_29 ? REG__2_cf_intrVec_2 : _GEN_3442; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3444 = 3'h3 == _T_29 ? REG__3_cf_intrVec_2 : _GEN_3443; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3445 = 3'h4 == _T_29 ? REG__4_cf_intrVec_2 : _GEN_3444; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3446 = 3'h5 == _T_29 ? REG__5_cf_intrVec_2 : _GEN_3445; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3447 = 3'h6 == _T_29 ? REG__6_cf_intrVec_2 : _GEN_3446; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3450 = 3'h1 == _T_29 ? REG__1_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3451 = 3'h2 == _T_29 ? REG__2_cf_intrVec_3 : _GEN_3450; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3452 = 3'h3 == _T_29 ? REG__3_cf_intrVec_3 : _GEN_3451; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3453 = 3'h4 == _T_29 ? REG__4_cf_intrVec_3 : _GEN_3452; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3454 = 3'h5 == _T_29 ? REG__5_cf_intrVec_3 : _GEN_3453; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3455 = 3'h6 == _T_29 ? REG__6_cf_intrVec_3 : _GEN_3454; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3458 = 3'h1 == _T_29 ? REG__1_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3459 = 3'h2 == _T_29 ? REG__2_cf_intrVec_4 : _GEN_3458; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3460 = 3'h3 == _T_29 ? REG__3_cf_intrVec_4 : _GEN_3459; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3461 = 3'h4 == _T_29 ? REG__4_cf_intrVec_4 : _GEN_3460; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3462 = 3'h5 == _T_29 ? REG__5_cf_intrVec_4 : _GEN_3461; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3463 = 3'h6 == _T_29 ? REG__6_cf_intrVec_4 : _GEN_3462; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3466 = 3'h1 == _T_29 ? REG__1_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3467 = 3'h2 == _T_29 ? REG__2_cf_intrVec_5 : _GEN_3466; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3468 = 3'h3 == _T_29 ? REG__3_cf_intrVec_5 : _GEN_3467; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3469 = 3'h4 == _T_29 ? REG__4_cf_intrVec_5 : _GEN_3468; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3470 = 3'h5 == _T_29 ? REG__5_cf_intrVec_5 : _GEN_3469; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3471 = 3'h6 == _T_29 ? REG__6_cf_intrVec_5 : _GEN_3470; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3474 = 3'h1 == _T_29 ? REG__1_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3475 = 3'h2 == _T_29 ? REG__2_cf_intrVec_6 : _GEN_3474; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3476 = 3'h3 == _T_29 ? REG__3_cf_intrVec_6 : _GEN_3475; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3477 = 3'h4 == _T_29 ? REG__4_cf_intrVec_6 : _GEN_3476; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3478 = 3'h5 == _T_29 ? REG__5_cf_intrVec_6 : _GEN_3477; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3479 = 3'h6 == _T_29 ? REG__6_cf_intrVec_6 : _GEN_3478; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3482 = 3'h1 == _T_29 ? REG__1_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3483 = 3'h2 == _T_29 ? REG__2_cf_intrVec_7 : _GEN_3482; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3484 = 3'h3 == _T_29 ? REG__3_cf_intrVec_7 : _GEN_3483; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3485 = 3'h4 == _T_29 ? REG__4_cf_intrVec_7 : _GEN_3484; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3486 = 3'h5 == _T_29 ? REG__5_cf_intrVec_7 : _GEN_3485; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3487 = 3'h6 == _T_29 ? REG__6_cf_intrVec_7 : _GEN_3486; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3490 = 3'h1 == _T_29 ? REG__1_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3491 = 3'h2 == _T_29 ? REG__2_cf_intrVec_8 : _GEN_3490; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3492 = 3'h3 == _T_29 ? REG__3_cf_intrVec_8 : _GEN_3491; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3493 = 3'h4 == _T_29 ? REG__4_cf_intrVec_8 : _GEN_3492; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3494 = 3'h5 == _T_29 ? REG__5_cf_intrVec_8 : _GEN_3493; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3495 = 3'h6 == _T_29 ? REG__6_cf_intrVec_8 : _GEN_3494; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3498 = 3'h1 == _T_29 ? REG__1_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3499 = 3'h2 == _T_29 ? REG__2_cf_intrVec_9 : _GEN_3498; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3500 = 3'h3 == _T_29 ? REG__3_cf_intrVec_9 : _GEN_3499; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3501 = 3'h4 == _T_29 ? REG__4_cf_intrVec_9 : _GEN_3500; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3502 = 3'h5 == _T_29 ? REG__5_cf_intrVec_9 : _GEN_3501; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3503 = 3'h6 == _T_29 ? REG__6_cf_intrVec_9 : _GEN_3502; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3506 = 3'h1 == _T_29 ? REG__1_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3507 = 3'h2 == _T_29 ? REG__2_cf_intrVec_10 : _GEN_3506; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3508 = 3'h3 == _T_29 ? REG__3_cf_intrVec_10 : _GEN_3507; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3509 = 3'h4 == _T_29 ? REG__4_cf_intrVec_10 : _GEN_3508; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3510 = 3'h5 == _T_29 ? REG__5_cf_intrVec_10 : _GEN_3509; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3511 = 3'h6 == _T_29 ? REG__6_cf_intrVec_10 : _GEN_3510; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3514 = 3'h1 == _T_29 ? REG__1_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3515 = 3'h2 == _T_29 ? REG__2_cf_intrVec_11 : _GEN_3514; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3516 = 3'h3 == _T_29 ? REG__3_cf_intrVec_11 : _GEN_3515; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3517 = 3'h4 == _T_29 ? REG__4_cf_intrVec_11 : _GEN_3516; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3518 = 3'h5 == _T_29 ? REG__5_cf_intrVec_11 : _GEN_3517; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3519 = 3'h6 == _T_29 ? REG__6_cf_intrVec_11 : _GEN_3518; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3530 = 3'h1 == _T_29 ? REG__1_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3531 = 3'h2 == _T_29 ? REG__2_cf_exceptionVec_1 : _GEN_3530; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3532 = 3'h3 == _T_29 ? REG__3_cf_exceptionVec_1 : _GEN_3531; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3533 = 3'h4 == _T_29 ? REG__4_cf_exceptionVec_1 : _GEN_3532; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3534 = 3'h5 == _T_29 ? REG__5_cf_exceptionVec_1 : _GEN_3533; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3535 = 3'h6 == _T_29 ? REG__6_cf_exceptionVec_1 : _GEN_3534; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3538 = 3'h1 == _T_29 ? REG__1_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3539 = 3'h2 == _T_29 ? REG__2_cf_exceptionVec_2 : _GEN_3538; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3540 = 3'h3 == _T_29 ? REG__3_cf_exceptionVec_2 : _GEN_3539; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3541 = 3'h4 == _T_29 ? REG__4_cf_exceptionVec_2 : _GEN_3540; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3542 = 3'h5 == _T_29 ? REG__5_cf_exceptionVec_2 : _GEN_3541; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3543 = 3'h6 == _T_29 ? REG__6_cf_exceptionVec_2 : _GEN_3542; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3618 = 3'h1 == _T_29 ? REG__1_cf_exceptionVec_12 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3619 = 3'h2 == _T_29 ? REG__2_cf_exceptionVec_12 : _GEN_3618; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3620 = 3'h3 == _T_29 ? REG__3_cf_exceptionVec_12 : _GEN_3619; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3621 = 3'h4 == _T_29 ? REG__4_cf_exceptionVec_12 : _GEN_3620; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3622 = 3'h5 == _T_29 ? REG__5_cf_exceptionVec_12 : _GEN_3621; // @[PipelineVector.scala 60:{15,15}]
  wire  _GEN_3623 = 3'h6 == _T_29 ? REG__6_cf_exceptionVec_12 : _GEN_3622; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3674 = 3'h1 == _T_29 ? REG__1_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3675 = 3'h2 == _T_29 ? REG__2_cf_pnpc : _GEN_3674; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3676 = 3'h3 == _T_29 ? REG__3_cf_pnpc : _GEN_3675; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3677 = 3'h4 == _T_29 ? REG__4_cf_pnpc : _GEN_3676; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3678 = 3'h5 == _T_29 ? REG__5_cf_pnpc : _GEN_3677; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3679 = 3'h6 == _T_29 ? REG__6_cf_pnpc : _GEN_3678; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3682 = 3'h1 == _T_29 ? REG__1_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3683 = 3'h2 == _T_29 ? REG__2_cf_pc : _GEN_3682; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3684 = 3'h3 == _T_29 ? REG__3_cf_pc : _GEN_3683; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3685 = 3'h4 == _T_29 ? REG__4_cf_pc : _GEN_3684; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3686 = 3'h5 == _T_29 ? REG__5_cf_pc : _GEN_3685; // @[PipelineVector.scala 60:{15,15}]
  wire [38:0] _GEN_3687 = 3'h6 == _T_29 ? REG__6_cf_pc : _GEN_3686; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3690 = 3'h1 == _T_29 ? REG__1_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3691 = 3'h2 == _T_29 ? REG__2_cf_instr : _GEN_3690; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3692 = 3'h3 == _T_29 ? REG__3_cf_instr : _GEN_3691; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3693 = 3'h4 == _T_29 ? REG__4_cf_instr : _GEN_3692; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3694 = 3'h5 == _T_29 ? REG__5_cf_instr : _GEN_3693; // @[PipelineVector.scala 60:{15,15}]
  wire [63:0] _GEN_3695 = 3'h6 == _T_29 ? REG__6_cf_instr : _GEN_3694; // @[PipelineVector.scala 60:{15,15}]
  wire  _T_32 = backend_io_in_0_ready & backend_io_in_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = backend_io_in_1_ready & backend_io_in_1_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_34 = _T_32 + _T_33; // @[PipelineVector.scala 64:44]
  wire  _T_35 = _T_34 > 2'h0; // @[PipelineVector.scala 65:35]
  wire [2:0] _GEN_3717 = {{1'd0}, _T_34}; // @[PipelineVector.scala 67:42]
  wire [2:0] _T_37 = REG_2 + _GEN_3717; // @[PipelineVector.scala 67:42]
  Frontend_inorder frontend ( // @[NutCore.scala 106:24]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(frontend_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_runahead_checkpoint_id(frontend_io_out_0_bits_cf_runahead_checkpoint_id),
    .io_out_0_bits_cf_instrType(frontend_io_out_0_bits_cf_instrType),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_funct3(frontend_io_out_0_bits_ctrl_funct3),
    .io_out_0_bits_ctrl_func24(frontend_io_out_0_bits_ctrl_func24),
    .io_out_0_bits_ctrl_func23(frontend_io_out_0_bits_ctrl_func23),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfSrc3(frontend_io_out_0_bits_ctrl_rfSrc3),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isMou(frontend_io_out_0_bits_ctrl_isMou),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .io_ipf(frontend_io_ipf),
    .flushICache(frontend_flushICache),
    .bpuUpdateReq_valid(frontend_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(frontend_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(frontend_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(frontend_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(frontend_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(frontend_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(frontend_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(frontend_bpuUpdateReq_isRVC),
    .vmEnable(frontend_vmEnable),
    .intrVec(frontend_intrVec),
    .flushTLB(frontend_flushTLB)
  );
  new_Backend_inorder backend ( // @[NutCore.scala 150:25]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_in_0_ready(backend_io_in_0_ready),
    .io_in_0_valid(backend_io_in_0_valid),
    .io_in_0_bits_cf_instr(backend_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(backend_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(backend_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(backend_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(backend_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(backend_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(backend_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(backend_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(backend_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(backend_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(backend_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(backend_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(backend_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(backend_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(backend_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(backend_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(backend_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(backend_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(backend_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(backend_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_cf_runahead_checkpoint_id(backend_io_in_0_bits_cf_runahead_checkpoint_id),
    .io_in_0_bits_cf_instrType(backend_io_in_0_bits_cf_instrType),
    .io_in_0_bits_ctrl_src1Type(backend_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(backend_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(backend_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(backend_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_funct3(backend_io_in_0_bits_ctrl_funct3),
    .io_in_0_bits_ctrl_func24(backend_io_in_0_bits_ctrl_func24),
    .io_in_0_bits_ctrl_func23(backend_io_in_0_bits_ctrl_func23),
    .io_in_0_bits_ctrl_rfSrc1(backend_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(backend_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfSrc3(backend_io_in_0_bits_ctrl_rfSrc3),
    .io_in_0_bits_ctrl_rfWen(backend_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(backend_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isMou(backend_io_in_0_bits_ctrl_isMou),
    .io_in_0_bits_data_imm(backend_io_in_0_bits_data_imm),
    .io_in_1_ready(backend_io_in_1_ready),
    .io_in_1_valid(backend_io_in_1_valid),
    .io_in_1_bits_cf_instr(backend_io_in_1_bits_cf_instr),
    .io_in_1_bits_cf_pc(backend_io_in_1_bits_cf_pc),
    .io_in_1_bits_cf_pnpc(backend_io_in_1_bits_cf_pnpc),
    .io_in_1_bits_cf_exceptionVec_1(backend_io_in_1_bits_cf_exceptionVec_1),
    .io_in_1_bits_cf_exceptionVec_2(backend_io_in_1_bits_cf_exceptionVec_2),
    .io_in_1_bits_cf_exceptionVec_12(backend_io_in_1_bits_cf_exceptionVec_12),
    .io_in_1_bits_cf_intrVec_0(backend_io_in_1_bits_cf_intrVec_0),
    .io_in_1_bits_cf_intrVec_1(backend_io_in_1_bits_cf_intrVec_1),
    .io_in_1_bits_cf_intrVec_2(backend_io_in_1_bits_cf_intrVec_2),
    .io_in_1_bits_cf_intrVec_3(backend_io_in_1_bits_cf_intrVec_3),
    .io_in_1_bits_cf_intrVec_4(backend_io_in_1_bits_cf_intrVec_4),
    .io_in_1_bits_cf_intrVec_5(backend_io_in_1_bits_cf_intrVec_5),
    .io_in_1_bits_cf_intrVec_6(backend_io_in_1_bits_cf_intrVec_6),
    .io_in_1_bits_cf_intrVec_7(backend_io_in_1_bits_cf_intrVec_7),
    .io_in_1_bits_cf_intrVec_8(backend_io_in_1_bits_cf_intrVec_8),
    .io_in_1_bits_cf_intrVec_9(backend_io_in_1_bits_cf_intrVec_9),
    .io_in_1_bits_cf_intrVec_10(backend_io_in_1_bits_cf_intrVec_10),
    .io_in_1_bits_cf_intrVec_11(backend_io_in_1_bits_cf_intrVec_11),
    .io_in_1_bits_cf_brIdx(backend_io_in_1_bits_cf_brIdx),
    .io_in_1_bits_cf_crossPageIPFFix(backend_io_in_1_bits_cf_crossPageIPFFix),
    .io_in_1_bits_cf_runahead_checkpoint_id(backend_io_in_1_bits_cf_runahead_checkpoint_id),
    .io_in_1_bits_cf_instrType(backend_io_in_1_bits_cf_instrType),
    .io_in_1_bits_ctrl_src1Type(backend_io_in_1_bits_ctrl_src1Type),
    .io_in_1_bits_ctrl_src2Type(backend_io_in_1_bits_ctrl_src2Type),
    .io_in_1_bits_ctrl_fuType(backend_io_in_1_bits_ctrl_fuType),
    .io_in_1_bits_ctrl_fuOpType(backend_io_in_1_bits_ctrl_fuOpType),
    .io_in_1_bits_ctrl_funct3(backend_io_in_1_bits_ctrl_funct3),
    .io_in_1_bits_ctrl_func24(backend_io_in_1_bits_ctrl_func24),
    .io_in_1_bits_ctrl_func23(backend_io_in_1_bits_ctrl_func23),
    .io_in_1_bits_ctrl_rfSrc1(backend_io_in_1_bits_ctrl_rfSrc1),
    .io_in_1_bits_ctrl_rfSrc2(backend_io_in_1_bits_ctrl_rfSrc2),
    .io_in_1_bits_ctrl_rfSrc3(backend_io_in_1_bits_ctrl_rfSrc3),
    .io_in_1_bits_ctrl_rfWen(backend_io_in_1_bits_ctrl_rfWen),
    .io_in_1_bits_ctrl_rfDest(backend_io_in_1_bits_ctrl_rfDest),
    .io_in_1_bits_ctrl_isMou(backend_io_in_1_bits_ctrl_isMou),
    .io_in_1_bits_data_imm(backend_io_in_1_bits_data_imm),
    .io_flush(backend_io_flush),
    .io_dmem_req_ready(backend_io_dmem_req_ready),
    .io_dmem_req_valid(backend_io_dmem_req_valid),
    .io_dmem_req_bits_addr(backend_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(backend_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(backend_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(backend_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(backend_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(backend_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(backend_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(backend_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(backend_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(backend_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(backend_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(backend_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(backend_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_addr(backend_io_memMMU_dmem_addr),
    .io_redirect_target(backend_io_redirect_target),
    .io_redirect_valid(backend_io_redirect_valid),
    ._T_408_0(backend__T_408_0),
    .flushICache(backend_flushICache),
    .perfCnts_2(backend_perfCnts_2),
    .io_in_0_bits_decode_cf_pc(backend_io_in_0_bits_decode_cf_pc),
    .satp(backend_satp),
    .bpuUpdateReq_valid(backend_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(backend_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(backend_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(backend_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(backend_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(backend_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(backend_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(backend_bpuUpdateReq_isRVC),
    .io_wb_rfDest_0(backend_io_wb_rfDest_0),
    .ismmio(backend_ismmio),
    .io_extra_mtip(backend_io_extra_mtip),
    .amoReq(backend_amoReq),
    .io_extra_meip_0(backend_io_extra_meip_0),
    .vmEnable(backend_vmEnable),
    .io_wb_rfWen_0(backend_io_wb_rfWen_0),
    .io_wb_WriteData_0(backend_io_wb_WriteData_0),
    .intrVec(backend_intrVec),
    ._T_407_0(backend__T_407_0),
    .io_extra_msip(backend_io_extra_msip),
    .flushTLB(backend_flushTLB),
    .io_in_0_valid_0(backend_io_in_0_valid_0)
  );
  SimpleBusCrossbarNto1 mmioXbar ( // @[NutCore.scala 158:26]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_0_req_ready(mmioXbar_io_in_0_req_ready),
    .io_in_0_req_valid(mmioXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(mmioXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(mmioXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(mmioXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(mmioXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(mmioXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(mmioXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(mmioXbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(mmioXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(mmioXbar_io_in_1_req_ready),
    .io_in_1_req_valid(mmioXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(mmioXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(mmioXbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(mmioXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(mmioXbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(mmioXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(mmioXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(mmioXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(mmioXbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(mmioXbar_io_out_req_ready),
    .io_out_req_valid(mmioXbar_io_out_req_valid),
    .io_out_req_bits_addr(mmioXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(mmioXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(mmioXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(mmioXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(mmioXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(mmioXbar_io_out_resp_ready),
    .io_out_resp_valid(mmioXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(mmioXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(mmioXbar_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 dmemXbar ( // @[NutCore.scala 159:26]
    .clock(dmemXbar_clock),
    .reset(dmemXbar_reset),
    .io_in_0_req_ready(dmemXbar_io_in_0_req_ready),
    .io_in_0_req_valid(dmemXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(dmemXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(dmemXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(dmemXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(dmemXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(dmemXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(dmemXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(dmemXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(dmemXbar_io_in_1_req_ready),
    .io_in_1_req_valid(dmemXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(dmemXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(dmemXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(dmemXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(dmemXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(dmemXbar_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(dmemXbar_io_in_2_req_ready),
    .io_in_2_req_valid(dmemXbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(dmemXbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(dmemXbar_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(dmemXbar_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(dmemXbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(dmemXbar_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(dmemXbar_io_in_3_req_ready),
    .io_in_3_req_valid(dmemXbar_io_in_3_req_valid),
    .io_in_3_req_bits_addr(dmemXbar_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(dmemXbar_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(dmemXbar_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(dmemXbar_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(dmemXbar_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(dmemXbar_io_in_3_resp_ready),
    .io_in_3_resp_valid(dmemXbar_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(dmemXbar_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(dmemXbar_io_in_3_resp_bits_rdata),
    .io_out_req_ready(dmemXbar_io_out_req_ready),
    .io_out_req_valid(dmemXbar_io_out_req_valid),
    .io_out_req_bits_addr(dmemXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(dmemXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(dmemXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dmemXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dmemXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(dmemXbar_io_out_resp_ready),
    .io_out_resp_valid(dmemXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(dmemXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dmemXbar_io_out_resp_bits_rdata)
  );
  SIMD_TLB itlb ( // @[EmbeddedTLB.scala 425:13]
    .clock(itlb_clock),
    .reset(itlb_reset),
    .io_in_req_ready(itlb_io_in_req_ready),
    .io_in_req_valid(itlb_io_in_req_valid),
    .io_in_req_bits_addr(itlb_io_in_req_bits_addr),
    .io_in_req_bits_user(itlb_io_in_req_bits_user),
    .io_in_resp_ready(itlb_io_in_resp_ready),
    .io_in_resp_valid(itlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(itlb_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(itlb_io_in_resp_bits_user),
    .io_out_req_ready(itlb_io_out_req_ready),
    .io_out_req_valid(itlb_io_out_req_valid),
    .io_out_req_bits_addr(itlb_io_out_req_bits_addr),
    .io_out_req_bits_size(itlb_io_out_req_bits_size),
    .io_out_req_bits_user(itlb_io_out_req_bits_user),
    .io_out_resp_ready(itlb_io_out_resp_ready),
    .io_out_resp_valid(itlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(itlb_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(itlb_io_out_resp_bits_user),
    .io_mem_req_ready(itlb_io_mem_req_ready),
    .io_mem_req_valid(itlb_io_mem_req_valid),
    .io_mem_req_bits_addr(itlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(itlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(itlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(itlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(itlb_io_mem_resp_bits_rdata),
    .io_flush(itlb_io_flush),
    .io_csrMMU_priviledgeMode(itlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_loadPF(itlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(itlb_io_csrMMU_storePF),
    .io_cacheEmpty(itlb_io_cacheEmpty),
    .io_ipf(itlb_io_ipf),
    .CSRSATP(itlb_CSRSATP),
    .MOUFlushTLB(itlb_MOUFlushTLB)
  );
  Cache Cache ( // @[Cache.scala 674:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_io_in_req_bits_size),
    .io_in_req_bits_user(Cache_io_in_req_bits_user),
    .io_in_resp_ready(Cache_io_in_resp_ready),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(Cache_io_in_resp_bits_user),
    .io_flush(Cache_io_flush),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(Cache_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_io_mmio_req_bits_size),
    .io_mmio_resp_valid(Cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_io_mmio_resp_bits_rdata),
    .io_empty(Cache_io_empty),
    .MOUFlushICache(Cache_MOUFlushICache)
  );
  SIMD_TLB_1 dtlb ( // @[EmbeddedTLB.scala 425:13]
    .clock(dtlb_clock),
    .reset(dtlb_reset),
    .io_in_req_ready(dtlb_io_in_req_ready),
    .io_in_req_valid(dtlb_io_in_req_valid),
    .io_in_req_bits_addr(dtlb_io_in_req_bits_addr),
    .io_in_req_bits_size(dtlb_io_in_req_bits_size),
    .io_in_req_bits_cmd(dtlb_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dtlb_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dtlb_io_in_req_bits_wdata),
    .io_in_resp_valid(dtlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(dtlb_io_in_resp_bits_rdata),
    .io_out_req_ready(dtlb_io_out_req_ready),
    .io_out_req_valid(dtlb_io_out_req_valid),
    .io_out_req_bits_addr(dtlb_io_out_req_bits_addr),
    .io_out_req_bits_size(dtlb_io_out_req_bits_size),
    .io_out_req_bits_cmd(dtlb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dtlb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dtlb_io_out_req_bits_wdata),
    .io_out_resp_valid(dtlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(dtlb_io_out_resp_bits_rdata),
    .io_mem_req_ready(dtlb_io_mem_req_ready),
    .io_mem_req_valid(dtlb_io_mem_req_valid),
    .io_mem_req_bits_addr(dtlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(dtlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(dtlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(dtlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(dtlb_io_mem_resp_bits_rdata),
    .io_flush(dtlb_io_flush),
    .io_csrMMU_priviledgeMode(dtlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(dtlb_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(dtlb_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(dtlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(dtlb_io_csrMMU_storePF),
    .io_csrMMU_addr(dtlb_io_csrMMU_addr),
    ._T_408_0(dtlb__T_408_0),
    .CSRSATP(dtlb_CSRSATP),
    .ismmio_0(dtlb_ismmio_0),
    .ISAMO(dtlb_ISAMO),
    .vmEnable_0(dtlb_vmEnable_0),
    ._T_407_0(dtlb__T_407_0),
    .MOUFlushTLB(dtlb_MOUFlushTLB)
  );
  Cache_1 Cache_1 ( // @[Cache.scala 674:35]
    .clock(Cache_1_clock),
    .reset(Cache_1_reset),
    .io_in_req_ready(Cache_1_io_in_req_ready),
    .io_in_req_valid(Cache_1_io_in_req_valid),
    .io_in_req_bits_addr(Cache_1_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_1_io_in_req_bits_wdata),
    .io_in_resp_ready(Cache_1_io_in_resp_ready),
    .io_in_resp_valid(Cache_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_1_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_1_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_1_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_1_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_1_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_1_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_1_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_1_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_1_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(Cache_1_io_out_coh_req_ready),
    .io_out_coh_req_valid(Cache_1_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(Cache_1_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(Cache_1_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_valid(Cache_1_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(Cache_1_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(Cache_1_io_out_coh_resp_bits_rdata),
    .io_mmio_req_ready(Cache_1_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_1_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_1_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_1_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(Cache_1_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(Cache_1_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(Cache_1_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(Cache_1_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_1_io_mmio_resp_bits_rdata)
  );
  assign io_imem_mem_req_valid = Cache_io_out_mem_req_valid; // @[NutCore.scala 163:13]
  assign io_imem_mem_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutCore.scala 163:13]
  assign io_imem_mem_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutCore.scala 163:13]
  assign io_imem_mem_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutCore.scala 163:13]
  assign io_dmem_mem_req_valid = Cache_1_io_out_mem_req_valid; // @[NutCore.scala 168:13]
  assign io_dmem_mem_req_bits_addr = Cache_1_io_out_mem_req_bits_addr; // @[NutCore.scala 168:13]
  assign io_dmem_mem_req_bits_cmd = Cache_1_io_out_mem_req_bits_cmd; // @[NutCore.scala 168:13]
  assign io_dmem_mem_req_bits_wdata = Cache_1_io_out_mem_req_bits_wdata; // @[NutCore.scala 168:13]
  assign io_dmem_coh_req_ready = Cache_1_io_out_coh_req_ready; // @[NutCore.scala 168:13]
  assign io_dmem_coh_resp_valid = Cache_1_io_out_coh_resp_valid; // @[NutCore.scala 168:13]
  assign io_dmem_coh_resp_bits_cmd = Cache_1_io_out_coh_resp_bits_cmd; // @[NutCore.scala 168:13]
  assign io_dmem_coh_resp_bits_rdata = Cache_1_io_out_coh_resp_bits_rdata; // @[NutCore.scala 168:13]
  assign io_mmio_req_valid = mmioXbar_io_out_req_valid; // @[NutCore.scala 177:13]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_req_bits_addr; // @[NutCore.scala 177:13]
  assign io_mmio_req_bits_size = mmioXbar_io_out_req_bits_size; // @[NutCore.scala 177:13]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_req_bits_cmd; // @[NutCore.scala 177:13]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_req_bits_wmask; // @[NutCore.scala 177:13]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_req_bits_wdata; // @[NutCore.scala 177:13]
  assign io_frontend_req_ready = dmemXbar_io_in_3_req_ready; // @[NutCore.scala 175:23]
  assign io_frontend_resp_valid = dmemXbar_io_in_3_resp_valid; // @[NutCore.scala 175:23]
  assign io_frontend_resp_bits_cmd = dmemXbar_io_in_3_resp_bits_cmd; // @[NutCore.scala 175:23]
  assign io_frontend_resp_bits_rdata = dmemXbar_io_in_3_resp_bits_rdata; // @[NutCore.scala 175:23]
  assign perfCnts_2 = backend_perfCnts_2;
  assign io_in_0_bits_decode_cf_pc = backend_io_in_0_bits_decode_cf_pc;
  assign io_wb_rfDest_0 = backend_io_wb_rfDest_0;
  assign io_wb_rfWen_0 = backend_io_wb_rfWen_0;
  assign io_wb_WriteData_0 = backend_io_wb_WriteData_0;
  assign io_in_0_valid_0 = backend_io_in_0_valid_0;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = itlb_io_in_req_ready; // @[EmbeddedTLB.scala 429:15]
  assign frontend_io_imem_resp_valid = itlb_io_in_resp_valid; // @[EmbeddedTLB.scala 429:15]
  assign frontend_io_imem_resp_bits_rdata = itlb_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 429:15]
  assign frontend_io_imem_resp_bits_user = itlb_io_in_resp_bits_user; // @[EmbeddedTLB.scala 429:15]
  assign frontend_io_out_0_ready = _T_9 | ~frontend_io_out_0_valid; // @[PipelineVector.scala 50:36]
  assign frontend_io_redirect_target = backend_io_redirect_target; // @[NutCore.scala 171:26]
  assign frontend_io_redirect_valid = backend_io_redirect_valid; // @[NutCore.scala 171:26]
  assign frontend_io_ipf = itlb_io_ipf; // @[NutCore.scala 162:21]
  assign frontend_flushICache = backend_flushICache;
  assign frontend_bpuUpdateReq_valid = backend_bpuUpdateReq_valid;
  assign frontend_bpuUpdateReq_pc = backend_bpuUpdateReq_pc;
  assign frontend_bpuUpdateReq_isMissPredict = backend_bpuUpdateReq_isMissPredict;
  assign frontend_bpuUpdateReq_actualTarget = backend_bpuUpdateReq_actualTarget;
  assign frontend_bpuUpdateReq_actualTaken = backend_bpuUpdateReq_actualTaken;
  assign frontend_bpuUpdateReq_fuOpType = backend_bpuUpdateReq_fuOpType;
  assign frontend_bpuUpdateReq_btbType = backend_bpuUpdateReq_btbType;
  assign frontend_bpuUpdateReq_isRVC = backend_bpuUpdateReq_isRVC;
  assign frontend_vmEnable = dtlb_vmEnable_0;
  assign frontend_intrVec = backend_intrVec;
  assign frontend_flushTLB = backend_flushTLB;
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_in_0_valid = REG_1 != REG_2; // @[PipelineVector.scala 56:34]
  assign backend_io_in_0_bits_cf_instr = 3'h7 == REG_2 ? REG__7_cf_instr : _GEN_3167; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pc = 3'h7 == REG_2 ? REG__7_cf_pc : _GEN_3159; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pnpc = 3'h7 == REG_2 ? REG__7_cf_pnpc : _GEN_3151; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_1 = 3'h7 == REG_2 ? REG__7_cf_exceptionVec_1 : _GEN_3007; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_2 = 3'h7 == REG_2 ? REG__7_cf_exceptionVec_2 : _GEN_3015; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_12 = 3'h7 == REG_2 ? REG__7_cf_exceptionVec_12 : _GEN_3095; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_0 = 3'h7 == REG_2 ? REG__7_cf_intrVec_0 : _GEN_2903; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_1 = 3'h7 == REG_2 ? REG__7_cf_intrVec_1 : _GEN_2911; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_2 = 3'h7 == REG_2 ? REG__7_cf_intrVec_2 : _GEN_2919; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_3 = 3'h7 == REG_2 ? REG__7_cf_intrVec_3 : _GEN_2927; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_4 = 3'h7 == REG_2 ? REG__7_cf_intrVec_4 : _GEN_2935; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_5 = 3'h7 == REG_2 ? REG__7_cf_intrVec_5 : _GEN_2943; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_6 = 3'h7 == REG_2 ? REG__7_cf_intrVec_6 : _GEN_2951; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_7 = 3'h7 == REG_2 ? REG__7_cf_intrVec_7 : _GEN_2959; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_8 = 3'h7 == REG_2 ? REG__7_cf_intrVec_8 : _GEN_2967; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_9 = 3'h7 == REG_2 ? REG__7_cf_intrVec_9 : _GEN_2975; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_10 = 3'h7 == REG_2 ? REG__7_cf_intrVec_10 : _GEN_2983; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_11 = 3'h7 == REG_2 ? REG__7_cf_intrVec_11 : _GEN_2991; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_brIdx = 3'h7 == REG_2 ? REG__7_cf_brIdx : _GEN_2895; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_crossPageIPFFix = 3'h7 == REG_2 ? REG__7_cf_crossPageIPFFix : _GEN_2879; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_runahead_checkpoint_id = 3'h7 == REG_2 ? REG__7_cf_runahead_checkpoint_id : _GEN_2871; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_instrType = 3'h7 == REG_2 ? REG__7_cf_instrType : _GEN_2855; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src1Type = 3'h7 == REG_2 ? REG__7_ctrl_src1Type : _GEN_2847; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src2Type = 3'h7 == REG_2 ? REG__7_ctrl_src2Type : _GEN_2839; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuType = 3'h7 == REG_2 ? REG__7_ctrl_fuType : _GEN_2831; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuOpType = 3'h7 == REG_2 ? REG__7_ctrl_fuOpType : _GEN_2823; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_funct3 = 3'h7 == REG_2 ? REG__7_ctrl_funct3 : _GEN_2815; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_func24 = 3'h7 == REG_2 ? REG__7_ctrl_func24 : _GEN_2807; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_func23 = 3'h7 == REG_2 ? REG__7_ctrl_func23 : _GEN_2799; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc1 = 3'h7 == REG_2 ? REG__7_ctrl_rfSrc1 : _GEN_2791; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc2 = 3'h7 == REG_2 ? REG__7_ctrl_rfSrc2 : _GEN_2783; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc3 = 3'h7 == REG_2 ? REG__7_ctrl_rfSrc3 : _GEN_2775; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfWen = 3'h7 == REG_2 ? REG__7_ctrl_rfWen : _GEN_2767; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfDest = 3'h7 == REG_2 ? REG__7_ctrl_rfDest : _GEN_2759; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_isMou = 3'h7 == REG_2 ? REG__7_ctrl_isMou : _GEN_2703; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_data_imm = 3'h7 == REG_2 ? REG__7_data_imm : _GEN_2671; // @[PipelineVector.scala 55:{15,15}]
  assign backend_io_in_1_valid = REG_1 != _T_29 & backend_io_in_0_valid; // @[PipelineVector.scala 61:54]
  assign backend_io_in_1_bits_cf_instr = 3'h7 == _T_29 ? REG__7_cf_instr : _GEN_3695; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_pc = 3'h7 == _T_29 ? REG__7_cf_pc : _GEN_3687; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_pnpc = 3'h7 == _T_29 ? REG__7_cf_pnpc : _GEN_3679; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_exceptionVec_1 = 3'h7 == _T_29 ? REG__7_cf_exceptionVec_1 : _GEN_3535; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_exceptionVec_2 = 3'h7 == _T_29 ? REG__7_cf_exceptionVec_2 : _GEN_3543; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_exceptionVec_12 = 3'h7 == _T_29 ? REG__7_cf_exceptionVec_12 : _GEN_3623; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_0 = 3'h7 == _T_29 ? REG__7_cf_intrVec_0 : _GEN_3431; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_1 = 3'h7 == _T_29 ? REG__7_cf_intrVec_1 : _GEN_3439; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_2 = 3'h7 == _T_29 ? REG__7_cf_intrVec_2 : _GEN_3447; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_3 = 3'h7 == _T_29 ? REG__7_cf_intrVec_3 : _GEN_3455; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_4 = 3'h7 == _T_29 ? REG__7_cf_intrVec_4 : _GEN_3463; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_5 = 3'h7 == _T_29 ? REG__7_cf_intrVec_5 : _GEN_3471; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_6 = 3'h7 == _T_29 ? REG__7_cf_intrVec_6 : _GEN_3479; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_7 = 3'h7 == _T_29 ? REG__7_cf_intrVec_7 : _GEN_3487; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_8 = 3'h7 == _T_29 ? REG__7_cf_intrVec_8 : _GEN_3495; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_9 = 3'h7 == _T_29 ? REG__7_cf_intrVec_9 : _GEN_3503; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_10 = 3'h7 == _T_29 ? REG__7_cf_intrVec_10 : _GEN_3511; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_intrVec_11 = 3'h7 == _T_29 ? REG__7_cf_intrVec_11 : _GEN_3519; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_brIdx = 3'h7 == _T_29 ? REG__7_cf_brIdx : _GEN_3423; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_crossPageIPFFix = 3'h7 == _T_29 ? REG__7_cf_crossPageIPFFix : _GEN_3407; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_runahead_checkpoint_id = 3'h7 == _T_29 ? REG__7_cf_runahead_checkpoint_id : _GEN_3399; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_cf_instrType = 3'h7 == _T_29 ? REG__7_cf_instrType : _GEN_3383; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_src1Type = 3'h7 == _T_29 ? REG__7_ctrl_src1Type : _GEN_3375; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_src2Type = 3'h7 == _T_29 ? REG__7_ctrl_src2Type : _GEN_3367; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_fuType = 3'h7 == _T_29 ? REG__7_ctrl_fuType : _GEN_3359; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_fuOpType = 3'h7 == _T_29 ? REG__7_ctrl_fuOpType : _GEN_3351; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_funct3 = 3'h7 == _T_29 ? REG__7_ctrl_funct3 : _GEN_3343; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_func24 = 3'h7 == _T_29 ? REG__7_ctrl_func24 : _GEN_3335; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_func23 = 3'h7 == _T_29 ? REG__7_ctrl_func23 : _GEN_3327; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_rfSrc1 = 3'h7 == _T_29 ? REG__7_ctrl_rfSrc1 : _GEN_3319; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_rfSrc2 = 3'h7 == _T_29 ? REG__7_ctrl_rfSrc2 : _GEN_3311; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_rfSrc3 = 3'h7 == _T_29 ? REG__7_ctrl_rfSrc3 : _GEN_3303; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_rfWen = 3'h7 == _T_29 ? REG__7_ctrl_rfWen : _GEN_3295; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_rfDest = 3'h7 == _T_29 ? REG__7_ctrl_rfDest : _GEN_3287; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_ctrl_isMou = 3'h7 == _T_29 ? REG__7_ctrl_isMou : _GEN_3231; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_in_1_bits_data_imm = 3'h7 == _T_29 ? REG__7_data_imm : _GEN_3199; // @[PipelineVector.scala 60:{15,15}]
  assign backend_io_flush = frontend_io_flushVec[3:2]; // @[NutCore.scala 172:45]
  assign backend_io_dmem_req_ready = dtlb_io_in_req_ready; // @[EmbeddedTLB.scala 429:15]
  assign backend_io_dmem_resp_valid = dtlb_io_in_resp_valid; // @[EmbeddedTLB.scala 429:15]
  assign backend_io_dmem_resp_bits_rdata = dtlb_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 429:15]
  assign backend_io_memMMU_dmem_loadPF = dtlb_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 432:19]
  assign backend_io_memMMU_dmem_storePF = dtlb_io_csrMMU_storePF; // @[EmbeddedTLB.scala 432:19]
  assign backend_io_memMMU_dmem_addr = dtlb_io_csrMMU_addr; // @[EmbeddedTLB.scala 432:19]
  assign backend__T_408_0 = dtlb__T_408_0;
  assign backend_ismmio = dtlb_ismmio_0;
  assign backend_io_extra_mtip = io_extra_mtip;
  assign backend_io_extra_meip_0 = io_extra_meip_0;
  assign backend_vmEnable = dtlb_vmEnable_0;
  assign backend__T_407_0 = dtlb__T_407_0;
  assign backend_io_extra_msip = io_extra_msip;
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_0_req_valid = Cache_io_mmio_req_valid; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_0_req_bits_addr = Cache_io_mmio_req_bits_addr; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_0_req_bits_size = Cache_io_mmio_req_bits_size; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_0_req_bits_cmd = 4'h0; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_0_req_bits_wmask = 8'h0; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_0_req_bits_wdata = 64'h0; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_1_req_valid = Cache_1_io_mmio_req_valid; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_1_req_bits_addr = Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_1_req_bits_size = Cache_1_io_mmio_req_bits_size; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_1_req_bits_cmd = Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_1_req_bits_wmask = Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 681:13]
  assign mmioXbar_io_in_1_req_bits_wdata = Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 681:13]
  assign mmioXbar_io_out_req_ready = io_mmio_req_ready; // @[NutCore.scala 177:13]
  assign mmioXbar_io_out_resp_valid = io_mmio_resp_valid; // @[NutCore.scala 177:13]
  assign mmioXbar_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[NutCore.scala 177:13]
  assign mmioXbar_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[NutCore.scala 177:13]
  assign dmemXbar_clock = clock;
  assign dmemXbar_reset = reset;
  assign dmemXbar_io_in_0_req_valid = dtlb_io_out_req_valid; // @[NutCore.scala 167:23]
  assign dmemXbar_io_in_0_req_bits_addr = dtlb_io_out_req_bits_addr; // @[NutCore.scala 167:23]
  assign dmemXbar_io_in_0_req_bits_size = dtlb_io_out_req_bits_size; // @[NutCore.scala 167:23]
  assign dmemXbar_io_in_0_req_bits_cmd = dtlb_io_out_req_bits_cmd; // @[NutCore.scala 167:23]
  assign dmemXbar_io_in_0_req_bits_wmask = dtlb_io_out_req_bits_wmask; // @[NutCore.scala 167:23]
  assign dmemXbar_io_in_0_req_bits_wdata = dtlb_io_out_req_bits_wdata; // @[NutCore.scala 167:23]
  assign dmemXbar_io_in_1_req_valid = itlb_io_mem_req_valid; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_1_req_bits_addr = itlb_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_1_req_bits_cmd = itlb_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_1_req_bits_wdata = itlb_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_2_req_valid = dtlb_io_mem_req_valid; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_2_req_bits_addr = dtlb_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_2_req_bits_cmd = dtlb_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_2_req_bits_wdata = dtlb_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 430:16]
  assign dmemXbar_io_in_3_req_valid = io_frontend_req_valid; // @[NutCore.scala 175:23]
  assign dmemXbar_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[NutCore.scala 175:23]
  assign dmemXbar_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[NutCore.scala 175:23]
  assign dmemXbar_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[NutCore.scala 175:23]
  assign dmemXbar_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[NutCore.scala 175:23]
  assign dmemXbar_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[NutCore.scala 175:23]
  assign dmemXbar_io_in_3_resp_ready = io_frontend_resp_ready; // @[NutCore.scala 175:23]
  assign dmemXbar_io_out_req_ready = Cache_1_io_in_req_ready; // @[Cache.scala 680:17]
  assign dmemXbar_io_out_resp_valid = Cache_1_io_in_resp_valid; // @[Cache.scala 680:17]
  assign dmemXbar_io_out_resp_bits_cmd = Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 680:17]
  assign dmemXbar_io_out_resp_bits_rdata = Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 680:17]
  assign itlb_clock = clock;
  assign itlb_reset = reset;
  assign itlb_io_in_req_valid = frontend_io_imem_req_valid; // @[EmbeddedTLB.scala 429:15]
  assign itlb_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[EmbeddedTLB.scala 429:15]
  assign itlb_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[EmbeddedTLB.scala 429:15]
  assign itlb_io_in_resp_ready = frontend_io_imem_resp_ready; // @[EmbeddedTLB.scala 429:15]
  assign itlb_io_out_req_ready = Cache_io_in_req_ready; // @[Cache.scala 680:17]
  assign itlb_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 680:17]
  assign itlb_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 680:17]
  assign itlb_io_out_resp_bits_user = Cache_io_in_resp_bits_user; // @[Cache.scala 680:17]
  assign itlb_io_mem_req_ready = dmemXbar_io_in_1_req_ready; // @[EmbeddedTLB.scala 430:16]
  assign itlb_io_mem_resp_valid = dmemXbar_io_in_1_resp_valid; // @[EmbeddedTLB.scala 430:16]
  assign itlb_io_mem_resp_bits_rdata = dmemXbar_io_in_1_resp_bits_rdata; // @[EmbeddedTLB.scala 430:16]
  assign itlb_io_flush = frontend_io_flushVec[0]; // @[NutCore.scala 161:104]
  assign itlb_io_csrMMU_priviledgeMode = backend_io_memMMU_imem_priviledgeMode; // @[EmbeddedTLB.scala 432:19]
  assign itlb_io_cacheEmpty = Cache_io_empty; // @[Cache.scala 682:11]
  assign itlb_CSRSATP = backend_satp;
  assign itlb_MOUFlushTLB = backend_flushTLB;
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = itlb_io_out_req_valid; // @[Cache.scala 680:17]
  assign Cache_io_in_req_bits_addr = itlb_io_out_req_bits_addr; // @[Cache.scala 680:17]
  assign Cache_io_in_req_bits_size = itlb_io_out_req_bits_size; // @[Cache.scala 680:17]
  assign Cache_io_in_req_bits_user = itlb_io_out_req_bits_user; // @[Cache.scala 680:17]
  assign Cache_io_in_resp_ready = itlb_io_out_resp_ready; // @[Cache.scala 680:17]
  assign Cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign Cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[NutCore.scala 163:13]
  assign Cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[NutCore.scala 163:13]
  assign Cache_io_out_mem_resp_bits_cmd = io_imem_mem_resp_bits_cmd; // @[NutCore.scala 163:13]
  assign Cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[NutCore.scala 163:13]
  assign Cache_io_mmio_req_ready = mmioXbar_io_in_0_req_ready; // @[Cache.scala 681:13]
  assign Cache_io_mmio_resp_valid = mmioXbar_io_in_0_resp_valid; // @[Cache.scala 681:13]
  assign Cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_0_resp_bits_rdata; // @[Cache.scala 681:13]
  assign Cache_MOUFlushICache = backend_flushICache;
  assign dtlb_clock = clock;
  assign dtlb_reset = reset;
  assign dtlb_io_in_req_valid = backend_io_dmem_req_valid; // @[EmbeddedTLB.scala 429:15]
  assign dtlb_io_in_req_bits_addr = backend_io_dmem_req_bits_addr; // @[EmbeddedTLB.scala 429:15]
  assign dtlb_io_in_req_bits_size = backend_io_dmem_req_bits_size; // @[EmbeddedTLB.scala 429:15]
  assign dtlb_io_in_req_bits_cmd = backend_io_dmem_req_bits_cmd; // @[EmbeddedTLB.scala 429:15]
  assign dtlb_io_in_req_bits_wmask = backend_io_dmem_req_bits_wmask; // @[EmbeddedTLB.scala 429:15]
  assign dtlb_io_in_req_bits_wdata = backend_io_dmem_req_bits_wdata; // @[EmbeddedTLB.scala 429:15]
  assign dtlb_io_out_req_ready = dmemXbar_io_in_0_req_ready; // @[NutCore.scala 167:23]
  assign dtlb_io_out_resp_valid = dmemXbar_io_in_0_resp_valid; // @[NutCore.scala 167:23]
  assign dtlb_io_out_resp_bits_rdata = dmemXbar_io_in_0_resp_bits_rdata; // @[NutCore.scala 167:23]
  assign dtlb_io_mem_req_ready = dmemXbar_io_in_2_req_ready; // @[EmbeddedTLB.scala 430:16]
  assign dtlb_io_mem_resp_valid = dmemXbar_io_in_2_resp_valid; // @[EmbeddedTLB.scala 430:16]
  assign dtlb_io_mem_resp_bits_rdata = dmemXbar_io_in_2_resp_bits_rdata; // @[EmbeddedTLB.scala 430:16]
  assign dtlb_io_flush = backend_io_flush[0]; // @[NutCore.scala 166:99]
  assign dtlb_io_csrMMU_priviledgeMode = backend_io_memMMU_dmem_priviledgeMode; // @[EmbeddedTLB.scala 432:19]
  assign dtlb_io_csrMMU_status_sum = backend_io_memMMU_dmem_status_sum; // @[EmbeddedTLB.scala 432:19]
  assign dtlb_io_csrMMU_status_mxr = backend_io_memMMU_dmem_status_mxr; // @[EmbeddedTLB.scala 432:19]
  assign dtlb_CSRSATP = backend_satp;
  assign dtlb_ISAMO = backend_amoReq;
  assign dtlb_MOUFlushTLB = backend_flushTLB;
  assign Cache_1_clock = clock;
  assign Cache_1_reset = reset;
  assign Cache_1_io_in_req_valid = dmemXbar_io_out_req_valid; // @[Cache.scala 680:17]
  assign Cache_1_io_in_req_bits_addr = dmemXbar_io_out_req_bits_addr; // @[Cache.scala 680:17]
  assign Cache_1_io_in_req_bits_size = dmemXbar_io_out_req_bits_size; // @[Cache.scala 680:17]
  assign Cache_1_io_in_req_bits_cmd = dmemXbar_io_out_req_bits_cmd; // @[Cache.scala 680:17]
  assign Cache_1_io_in_req_bits_wmask = dmemXbar_io_out_req_bits_wmask; // @[Cache.scala 680:17]
  assign Cache_1_io_in_req_bits_wdata = dmemXbar_io_out_req_bits_wdata; // @[Cache.scala 680:17]
  assign Cache_1_io_in_resp_ready = dmemXbar_io_out_resp_ready; // @[Cache.scala 680:17]
  assign Cache_1_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[NutCore.scala 168:13]
  assign Cache_1_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[NutCore.scala 168:13]
  assign Cache_1_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[NutCore.scala 168:13]
  assign Cache_1_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[NutCore.scala 168:13]
  assign Cache_1_io_out_coh_req_valid = io_dmem_coh_req_valid; // @[NutCore.scala 168:13]
  assign Cache_1_io_out_coh_req_bits_addr = io_dmem_coh_req_bits_addr; // @[NutCore.scala 168:13]
  assign Cache_1_io_out_coh_req_bits_wdata = io_dmem_coh_req_bits_wdata; // @[NutCore.scala 168:13]
  assign Cache_1_io_mmio_req_ready = mmioXbar_io_in_1_req_ready; // @[Cache.scala 681:13]
  assign Cache_1_io_mmio_resp_valid = mmioXbar_io_in_1_resp_valid; // @[Cache.scala 681:13]
  assign Cache_1_io_mmio_resp_bits_rdata = mmioXbar_io_in_1_resp_bits_rdata; // @[Cache.scala 681:13]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_instr <= _GEN_1048;
        end
      end else begin
        REG__0_cf_instr <= _GEN_1048;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_pc <= _GEN_1040;
        end
      end else begin
        REG__0_cf_pc <= _GEN_1040;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_pnpc <= _GEN_1032;
        end
      end else begin
        REG__0_cf_pnpc <= _GEN_1032;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_1 <= _GEN_888;
        end
      end else begin
        REG__0_cf_exceptionVec_1 <= _GEN_888;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_2 <= _GEN_896;
        end
      end else begin
        REG__0_cf_exceptionVec_2 <= _GEN_896;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_12 <= _GEN_976;
        end
      end else begin
        REG__0_cf_exceptionVec_12 <= _GEN_976;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_0 <= _GEN_784;
        end
      end else begin
        REG__0_cf_intrVec_0 <= _GEN_784;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_1 <= _GEN_792;
        end
      end else begin
        REG__0_cf_intrVec_1 <= _GEN_792;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_2 <= _GEN_800;
        end
      end else begin
        REG__0_cf_intrVec_2 <= _GEN_800;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_3 <= _GEN_808;
        end
      end else begin
        REG__0_cf_intrVec_3 <= _GEN_808;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_4 <= _GEN_816;
        end
      end else begin
        REG__0_cf_intrVec_4 <= _GEN_816;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_5 <= _GEN_824;
        end
      end else begin
        REG__0_cf_intrVec_5 <= _GEN_824;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_6 <= _GEN_832;
        end
      end else begin
        REG__0_cf_intrVec_6 <= _GEN_832;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_7 <= _GEN_840;
        end
      end else begin
        REG__0_cf_intrVec_7 <= _GEN_840;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_8 <= _GEN_848;
        end
      end else begin
        REG__0_cf_intrVec_8 <= _GEN_848;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_9 <= _GEN_856;
        end
      end else begin
        REG__0_cf_intrVec_9 <= _GEN_856;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_10 <= _GEN_864;
        end
      end else begin
        REG__0_cf_intrVec_10 <= _GEN_864;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_11 <= _GEN_872;
        end
      end else begin
        REG__0_cf_intrVec_11 <= _GEN_872;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_brIdx <= _GEN_776;
        end
      end else begin
        REG__0_cf_brIdx <= _GEN_776;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_crossPageIPFFix <= _GEN_760;
        end
      end else begin
        REG__0_cf_crossPageIPFFix <= _GEN_760;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_runahead_checkpoint_id <= _GEN_752;
        end
      end else begin
        REG__0_cf_runahead_checkpoint_id <= _GEN_752;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_instrType <= _GEN_736;
        end
      end else begin
        REG__0_cf_instrType <= _GEN_736;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__0_ctrl_src1Type <= 3'h0 == _T_20 | _GEN_728;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__0_ctrl_src1Type <= _GEN_200;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__0_ctrl_src2Type <= 3'h0 == _T_20 | _GEN_720;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__0_ctrl_src2Type <= _GEN_192;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_fuType <= _GEN_712;
        end
      end else begin
        REG__0_ctrl_fuType <= _GEN_712;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_fuOpType <= _GEN_704;
        end
      end else begin
        REG__0_ctrl_fuOpType <= _GEN_704;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_funct3 <= _GEN_696;
        end
      end else begin
        REG__0_ctrl_funct3 <= _GEN_696;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_func24 <= _GEN_688;
        end
      end else begin
        REG__0_ctrl_func24 <= _GEN_688;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_func23 <= _GEN_680;
        end
      end else begin
        REG__0_ctrl_func23 <= _GEN_680;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc1 <= _GEN_672;
        end
      end else begin
        REG__0_ctrl_rfSrc1 <= _GEN_672;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc2 <= _GEN_664;
        end
      end else begin
        REG__0_ctrl_rfSrc2 <= _GEN_664;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc3 <= _GEN_656;
        end
      end else begin
        REG__0_ctrl_rfSrc3 <= _GEN_656;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfWen <= _GEN_648;
        end
      end else begin
        REG__0_ctrl_rfWen <= _GEN_648;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfDest <= _GEN_640;
        end
      end else begin
        REG__0_ctrl_rfDest <= _GEN_640;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_isMou <= _GEN_584;
        end
      end else begin
        REG__0_ctrl_isMou <= _GEN_584;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_data_imm <= _GEN_552;
        end
      end else begin
        REG__0_data_imm <= _GEN_552;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_instr <= _GEN_1049;
        end
      end else begin
        REG__1_cf_instr <= _GEN_1049;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_pc <= _GEN_1041;
        end
      end else begin
        REG__1_cf_pc <= _GEN_1041;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_pnpc <= _GEN_1033;
        end
      end else begin
        REG__1_cf_pnpc <= _GEN_1033;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_1 <= _GEN_889;
        end
      end else begin
        REG__1_cf_exceptionVec_1 <= _GEN_889;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_2 <= _GEN_897;
        end
      end else begin
        REG__1_cf_exceptionVec_2 <= _GEN_897;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_12 <= _GEN_977;
        end
      end else begin
        REG__1_cf_exceptionVec_12 <= _GEN_977;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_0 <= _GEN_785;
        end
      end else begin
        REG__1_cf_intrVec_0 <= _GEN_785;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_1 <= _GEN_793;
        end
      end else begin
        REG__1_cf_intrVec_1 <= _GEN_793;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_2 <= _GEN_801;
        end
      end else begin
        REG__1_cf_intrVec_2 <= _GEN_801;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_3 <= _GEN_809;
        end
      end else begin
        REG__1_cf_intrVec_3 <= _GEN_809;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_4 <= _GEN_817;
        end
      end else begin
        REG__1_cf_intrVec_4 <= _GEN_817;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_5 <= _GEN_825;
        end
      end else begin
        REG__1_cf_intrVec_5 <= _GEN_825;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_6 <= _GEN_833;
        end
      end else begin
        REG__1_cf_intrVec_6 <= _GEN_833;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_7 <= _GEN_841;
        end
      end else begin
        REG__1_cf_intrVec_7 <= _GEN_841;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_8 <= _GEN_849;
        end
      end else begin
        REG__1_cf_intrVec_8 <= _GEN_849;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_9 <= _GEN_857;
        end
      end else begin
        REG__1_cf_intrVec_9 <= _GEN_857;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_10 <= _GEN_865;
        end
      end else begin
        REG__1_cf_intrVec_10 <= _GEN_865;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_11 <= _GEN_873;
        end
      end else begin
        REG__1_cf_intrVec_11 <= _GEN_873;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_brIdx <= _GEN_777;
        end
      end else begin
        REG__1_cf_brIdx <= _GEN_777;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_crossPageIPFFix <= _GEN_761;
        end
      end else begin
        REG__1_cf_crossPageIPFFix <= _GEN_761;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_runahead_checkpoint_id <= _GEN_753;
        end
      end else begin
        REG__1_cf_runahead_checkpoint_id <= _GEN_753;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_instrType <= _GEN_737;
        end
      end else begin
        REG__1_cf_instrType <= _GEN_737;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__1_ctrl_src1Type <= 3'h1 == _T_20 | _GEN_729;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__1_ctrl_src1Type <= _GEN_201;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__1_ctrl_src2Type <= 3'h1 == _T_20 | _GEN_721;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__1_ctrl_src2Type <= _GEN_193;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_fuType <= _GEN_713;
        end
      end else begin
        REG__1_ctrl_fuType <= _GEN_713;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_fuOpType <= _GEN_705;
        end
      end else begin
        REG__1_ctrl_fuOpType <= _GEN_705;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_funct3 <= _GEN_697;
        end
      end else begin
        REG__1_ctrl_funct3 <= _GEN_697;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_func24 <= _GEN_689;
        end
      end else begin
        REG__1_ctrl_func24 <= _GEN_689;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_func23 <= _GEN_681;
        end
      end else begin
        REG__1_ctrl_func23 <= _GEN_681;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc1 <= _GEN_673;
        end
      end else begin
        REG__1_ctrl_rfSrc1 <= _GEN_673;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc2 <= _GEN_665;
        end
      end else begin
        REG__1_ctrl_rfSrc2 <= _GEN_665;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc3 <= _GEN_657;
        end
      end else begin
        REG__1_ctrl_rfSrc3 <= _GEN_657;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfWen <= _GEN_649;
        end
      end else begin
        REG__1_ctrl_rfWen <= _GEN_649;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfDest <= _GEN_641;
        end
      end else begin
        REG__1_ctrl_rfDest <= _GEN_641;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_isMou <= _GEN_585;
        end
      end else begin
        REG__1_ctrl_isMou <= _GEN_585;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_data_imm <= _GEN_553;
        end
      end else begin
        REG__1_data_imm <= _GEN_553;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_instr <= _GEN_1050;
        end
      end else begin
        REG__2_cf_instr <= _GEN_1050;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_pc <= _GEN_1042;
        end
      end else begin
        REG__2_cf_pc <= _GEN_1042;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_pnpc <= _GEN_1034;
        end
      end else begin
        REG__2_cf_pnpc <= _GEN_1034;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_1 <= _GEN_890;
        end
      end else begin
        REG__2_cf_exceptionVec_1 <= _GEN_890;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_2 <= _GEN_898;
        end
      end else begin
        REG__2_cf_exceptionVec_2 <= _GEN_898;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_12 <= _GEN_978;
        end
      end else begin
        REG__2_cf_exceptionVec_12 <= _GEN_978;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_0 <= _GEN_786;
        end
      end else begin
        REG__2_cf_intrVec_0 <= _GEN_786;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_1 <= _GEN_794;
        end
      end else begin
        REG__2_cf_intrVec_1 <= _GEN_794;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_2 <= _GEN_802;
        end
      end else begin
        REG__2_cf_intrVec_2 <= _GEN_802;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_3 <= _GEN_810;
        end
      end else begin
        REG__2_cf_intrVec_3 <= _GEN_810;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_4 <= _GEN_818;
        end
      end else begin
        REG__2_cf_intrVec_4 <= _GEN_818;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_5 <= _GEN_826;
        end
      end else begin
        REG__2_cf_intrVec_5 <= _GEN_826;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_6 <= _GEN_834;
        end
      end else begin
        REG__2_cf_intrVec_6 <= _GEN_834;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_7 <= _GEN_842;
        end
      end else begin
        REG__2_cf_intrVec_7 <= _GEN_842;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_8 <= _GEN_850;
        end
      end else begin
        REG__2_cf_intrVec_8 <= _GEN_850;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_9 <= _GEN_858;
        end
      end else begin
        REG__2_cf_intrVec_9 <= _GEN_858;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_10 <= _GEN_866;
        end
      end else begin
        REG__2_cf_intrVec_10 <= _GEN_866;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_11 <= _GEN_874;
        end
      end else begin
        REG__2_cf_intrVec_11 <= _GEN_874;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_brIdx <= _GEN_778;
        end
      end else begin
        REG__2_cf_brIdx <= _GEN_778;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_crossPageIPFFix <= _GEN_762;
        end
      end else begin
        REG__2_cf_crossPageIPFFix <= _GEN_762;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_runahead_checkpoint_id <= _GEN_754;
        end
      end else begin
        REG__2_cf_runahead_checkpoint_id <= _GEN_754;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_instrType <= _GEN_738;
        end
      end else begin
        REG__2_cf_instrType <= _GEN_738;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__2_ctrl_src1Type <= 3'h2 == _T_20 | _GEN_730;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__2_ctrl_src1Type <= _GEN_202;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__2_ctrl_src2Type <= 3'h2 == _T_20 | _GEN_722;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__2_ctrl_src2Type <= _GEN_194;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_fuType <= _GEN_714;
        end
      end else begin
        REG__2_ctrl_fuType <= _GEN_714;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_fuOpType <= _GEN_706;
        end
      end else begin
        REG__2_ctrl_fuOpType <= _GEN_706;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_funct3 <= _GEN_698;
        end
      end else begin
        REG__2_ctrl_funct3 <= _GEN_698;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_func24 <= _GEN_690;
        end
      end else begin
        REG__2_ctrl_func24 <= _GEN_690;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_func23 <= _GEN_682;
        end
      end else begin
        REG__2_ctrl_func23 <= _GEN_682;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc1 <= _GEN_674;
        end
      end else begin
        REG__2_ctrl_rfSrc1 <= _GEN_674;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc2 <= _GEN_666;
        end
      end else begin
        REG__2_ctrl_rfSrc2 <= _GEN_666;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc3 <= _GEN_658;
        end
      end else begin
        REG__2_ctrl_rfSrc3 <= _GEN_658;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfWen <= _GEN_650;
        end
      end else begin
        REG__2_ctrl_rfWen <= _GEN_650;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfDest <= _GEN_642;
        end
      end else begin
        REG__2_ctrl_rfDest <= _GEN_642;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_isMou <= _GEN_586;
        end
      end else begin
        REG__2_ctrl_isMou <= _GEN_586;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_data_imm <= _GEN_554;
        end
      end else begin
        REG__2_data_imm <= _GEN_554;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_instr <= _GEN_1051;
        end
      end else begin
        REG__3_cf_instr <= _GEN_1051;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_pc <= _GEN_1043;
        end
      end else begin
        REG__3_cf_pc <= _GEN_1043;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_pnpc <= _GEN_1035;
        end
      end else begin
        REG__3_cf_pnpc <= _GEN_1035;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_1 <= _GEN_891;
        end
      end else begin
        REG__3_cf_exceptionVec_1 <= _GEN_891;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_2 <= _GEN_899;
        end
      end else begin
        REG__3_cf_exceptionVec_2 <= _GEN_899;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_12 <= _GEN_979;
        end
      end else begin
        REG__3_cf_exceptionVec_12 <= _GEN_979;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_0 <= _GEN_787;
        end
      end else begin
        REG__3_cf_intrVec_0 <= _GEN_787;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_1 <= _GEN_795;
        end
      end else begin
        REG__3_cf_intrVec_1 <= _GEN_795;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_2 <= _GEN_803;
        end
      end else begin
        REG__3_cf_intrVec_2 <= _GEN_803;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_3 <= _GEN_811;
        end
      end else begin
        REG__3_cf_intrVec_3 <= _GEN_811;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_4 <= _GEN_819;
        end
      end else begin
        REG__3_cf_intrVec_4 <= _GEN_819;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_5 <= _GEN_827;
        end
      end else begin
        REG__3_cf_intrVec_5 <= _GEN_827;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_6 <= _GEN_835;
        end
      end else begin
        REG__3_cf_intrVec_6 <= _GEN_835;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_7 <= _GEN_843;
        end
      end else begin
        REG__3_cf_intrVec_7 <= _GEN_843;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_8 <= _GEN_851;
        end
      end else begin
        REG__3_cf_intrVec_8 <= _GEN_851;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_9 <= _GEN_859;
        end
      end else begin
        REG__3_cf_intrVec_9 <= _GEN_859;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_10 <= _GEN_867;
        end
      end else begin
        REG__3_cf_intrVec_10 <= _GEN_867;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_11 <= _GEN_875;
        end
      end else begin
        REG__3_cf_intrVec_11 <= _GEN_875;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_brIdx <= _GEN_779;
        end
      end else begin
        REG__3_cf_brIdx <= _GEN_779;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_crossPageIPFFix <= _GEN_763;
        end
      end else begin
        REG__3_cf_crossPageIPFFix <= _GEN_763;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_runahead_checkpoint_id <= _GEN_755;
        end
      end else begin
        REG__3_cf_runahead_checkpoint_id <= _GEN_755;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_instrType <= _GEN_739;
        end
      end else begin
        REG__3_cf_instrType <= _GEN_739;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__3_ctrl_src1Type <= 3'h3 == _T_20 | _GEN_731;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__3_ctrl_src1Type <= _GEN_203;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__3_ctrl_src2Type <= 3'h3 == _T_20 | _GEN_723;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__3_ctrl_src2Type <= _GEN_195;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_fuType <= _GEN_715;
        end
      end else begin
        REG__3_ctrl_fuType <= _GEN_715;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_fuOpType <= _GEN_707;
        end
      end else begin
        REG__3_ctrl_fuOpType <= _GEN_707;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_funct3 <= _GEN_699;
        end
      end else begin
        REG__3_ctrl_funct3 <= _GEN_699;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_func24 <= _GEN_691;
        end
      end else begin
        REG__3_ctrl_func24 <= _GEN_691;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_func23 <= _GEN_683;
        end
      end else begin
        REG__3_ctrl_func23 <= _GEN_683;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc1 <= _GEN_675;
        end
      end else begin
        REG__3_ctrl_rfSrc1 <= _GEN_675;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc2 <= _GEN_667;
        end
      end else begin
        REG__3_ctrl_rfSrc2 <= _GEN_667;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc3 <= _GEN_659;
        end
      end else begin
        REG__3_ctrl_rfSrc3 <= _GEN_659;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfWen <= _GEN_651;
        end
      end else begin
        REG__3_ctrl_rfWen <= _GEN_651;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfDest <= _GEN_643;
        end
      end else begin
        REG__3_ctrl_rfDest <= _GEN_643;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_isMou <= _GEN_587;
        end
      end else begin
        REG__3_ctrl_isMou <= _GEN_587;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_data_imm <= _GEN_555;
        end
      end else begin
        REG__3_data_imm <= _GEN_555;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_instr <= _GEN_1052;
        end
      end else begin
        REG__4_cf_instr <= _GEN_1052;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_pc <= _GEN_1044;
        end
      end else begin
        REG__4_cf_pc <= _GEN_1044;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_pnpc <= _GEN_1036;
        end
      end else begin
        REG__4_cf_pnpc <= _GEN_1036;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_exceptionVec_1 <= _GEN_892;
        end
      end else begin
        REG__4_cf_exceptionVec_1 <= _GEN_892;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_exceptionVec_2 <= _GEN_900;
        end
      end else begin
        REG__4_cf_exceptionVec_2 <= _GEN_900;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_exceptionVec_12 <= _GEN_980;
        end
      end else begin
        REG__4_cf_exceptionVec_12 <= _GEN_980;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_0 <= _GEN_788;
        end
      end else begin
        REG__4_cf_intrVec_0 <= _GEN_788;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_1 <= _GEN_796;
        end
      end else begin
        REG__4_cf_intrVec_1 <= _GEN_796;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_2 <= _GEN_804;
        end
      end else begin
        REG__4_cf_intrVec_2 <= _GEN_804;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_3 <= _GEN_812;
        end
      end else begin
        REG__4_cf_intrVec_3 <= _GEN_812;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_4 <= _GEN_820;
        end
      end else begin
        REG__4_cf_intrVec_4 <= _GEN_820;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_5 <= _GEN_828;
        end
      end else begin
        REG__4_cf_intrVec_5 <= _GEN_828;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_6 <= _GEN_836;
        end
      end else begin
        REG__4_cf_intrVec_6 <= _GEN_836;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_7 <= _GEN_844;
        end
      end else begin
        REG__4_cf_intrVec_7 <= _GEN_844;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_8 <= _GEN_852;
        end
      end else begin
        REG__4_cf_intrVec_8 <= _GEN_852;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_9 <= _GEN_860;
        end
      end else begin
        REG__4_cf_intrVec_9 <= _GEN_860;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_10 <= _GEN_868;
        end
      end else begin
        REG__4_cf_intrVec_10 <= _GEN_868;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_intrVec_11 <= _GEN_876;
        end
      end else begin
        REG__4_cf_intrVec_11 <= _GEN_876;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_brIdx <= _GEN_780;
        end
      end else begin
        REG__4_cf_brIdx <= _GEN_780;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_crossPageIPFFix <= _GEN_764;
        end
      end else begin
        REG__4_cf_crossPageIPFFix <= _GEN_764;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_runahead_checkpoint_id <= _GEN_756;
        end
      end else begin
        REG__4_cf_runahead_checkpoint_id <= _GEN_756;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_cf_instrType <= _GEN_740;
        end
      end else begin
        REG__4_cf_instrType <= _GEN_740;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__4_ctrl_src1Type <= 3'h4 == _T_20 | _GEN_732;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__4_ctrl_src1Type <= _GEN_204;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__4_ctrl_src2Type <= 3'h4 == _T_20 | _GEN_724;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__4_ctrl_src2Type <= _GEN_196;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_fuType <= _GEN_716;
        end
      end else begin
        REG__4_ctrl_fuType <= _GEN_716;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_fuOpType <= _GEN_708;
        end
      end else begin
        REG__4_ctrl_fuOpType <= _GEN_708;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_funct3 <= _GEN_700;
        end
      end else begin
        REG__4_ctrl_funct3 <= _GEN_700;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_func24 <= _GEN_692;
        end
      end else begin
        REG__4_ctrl_func24 <= _GEN_692;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_func23 <= _GEN_684;
        end
      end else begin
        REG__4_ctrl_func23 <= _GEN_684;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_rfSrc1 <= _GEN_676;
        end
      end else begin
        REG__4_ctrl_rfSrc1 <= _GEN_676;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_rfSrc2 <= _GEN_668;
        end
      end else begin
        REG__4_ctrl_rfSrc2 <= _GEN_668;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_rfSrc3 <= _GEN_660;
        end
      end else begin
        REG__4_ctrl_rfSrc3 <= _GEN_660;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_rfWen <= _GEN_652;
        end
      end else begin
        REG__4_ctrl_rfWen <= _GEN_652;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_rfDest <= _GEN_644;
        end
      end else begin
        REG__4_ctrl_rfDest <= _GEN_644;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_ctrl_isMou <= _GEN_588;
        end
      end else begin
        REG__4_ctrl_isMou <= _GEN_588;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__4_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h4 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__4_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__4_data_imm <= _GEN_556;
        end
      end else begin
        REG__4_data_imm <= _GEN_556;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_instr <= _GEN_1053;
        end
      end else begin
        REG__5_cf_instr <= _GEN_1053;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_pc <= _GEN_1045;
        end
      end else begin
        REG__5_cf_pc <= _GEN_1045;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_pnpc <= _GEN_1037;
        end
      end else begin
        REG__5_cf_pnpc <= _GEN_1037;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_exceptionVec_1 <= _GEN_893;
        end
      end else begin
        REG__5_cf_exceptionVec_1 <= _GEN_893;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_exceptionVec_2 <= _GEN_901;
        end
      end else begin
        REG__5_cf_exceptionVec_2 <= _GEN_901;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_exceptionVec_12 <= _GEN_981;
        end
      end else begin
        REG__5_cf_exceptionVec_12 <= _GEN_981;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_0 <= _GEN_789;
        end
      end else begin
        REG__5_cf_intrVec_0 <= _GEN_789;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_1 <= _GEN_797;
        end
      end else begin
        REG__5_cf_intrVec_1 <= _GEN_797;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_2 <= _GEN_805;
        end
      end else begin
        REG__5_cf_intrVec_2 <= _GEN_805;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_3 <= _GEN_813;
        end
      end else begin
        REG__5_cf_intrVec_3 <= _GEN_813;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_4 <= _GEN_821;
        end
      end else begin
        REG__5_cf_intrVec_4 <= _GEN_821;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_5 <= _GEN_829;
        end
      end else begin
        REG__5_cf_intrVec_5 <= _GEN_829;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_6 <= _GEN_837;
        end
      end else begin
        REG__5_cf_intrVec_6 <= _GEN_837;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_7 <= _GEN_845;
        end
      end else begin
        REG__5_cf_intrVec_7 <= _GEN_845;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_8 <= _GEN_853;
        end
      end else begin
        REG__5_cf_intrVec_8 <= _GEN_853;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_9 <= _GEN_861;
        end
      end else begin
        REG__5_cf_intrVec_9 <= _GEN_861;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_10 <= _GEN_869;
        end
      end else begin
        REG__5_cf_intrVec_10 <= _GEN_869;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_intrVec_11 <= _GEN_877;
        end
      end else begin
        REG__5_cf_intrVec_11 <= _GEN_877;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_brIdx <= _GEN_781;
        end
      end else begin
        REG__5_cf_brIdx <= _GEN_781;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_crossPageIPFFix <= _GEN_765;
        end
      end else begin
        REG__5_cf_crossPageIPFFix <= _GEN_765;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_runahead_checkpoint_id <= _GEN_757;
        end
      end else begin
        REG__5_cf_runahead_checkpoint_id <= _GEN_757;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_cf_instrType <= _GEN_741;
        end
      end else begin
        REG__5_cf_instrType <= _GEN_741;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__5_ctrl_src1Type <= 3'h5 == _T_20 | _GEN_733;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__5_ctrl_src1Type <= _GEN_205;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__5_ctrl_src2Type <= 3'h5 == _T_20 | _GEN_725;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__5_ctrl_src2Type <= _GEN_197;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_fuType <= _GEN_717;
        end
      end else begin
        REG__5_ctrl_fuType <= _GEN_717;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_fuOpType <= _GEN_709;
        end
      end else begin
        REG__5_ctrl_fuOpType <= _GEN_709;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_funct3 <= _GEN_701;
        end
      end else begin
        REG__5_ctrl_funct3 <= _GEN_701;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_func24 <= _GEN_693;
        end
      end else begin
        REG__5_ctrl_func24 <= _GEN_693;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_func23 <= _GEN_685;
        end
      end else begin
        REG__5_ctrl_func23 <= _GEN_685;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_rfSrc1 <= _GEN_677;
        end
      end else begin
        REG__5_ctrl_rfSrc1 <= _GEN_677;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_rfSrc2 <= _GEN_669;
        end
      end else begin
        REG__5_ctrl_rfSrc2 <= _GEN_669;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_rfSrc3 <= _GEN_661;
        end
      end else begin
        REG__5_ctrl_rfSrc3 <= _GEN_661;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_rfWen <= _GEN_653;
        end
      end else begin
        REG__5_ctrl_rfWen <= _GEN_653;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_rfDest <= _GEN_645;
        end
      end else begin
        REG__5_ctrl_rfDest <= _GEN_645;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_ctrl_isMou <= _GEN_589;
        end
      end else begin
        REG__5_ctrl_isMou <= _GEN_589;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__5_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h5 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__5_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__5_data_imm <= _GEN_557;
        end
      end else begin
        REG__5_data_imm <= _GEN_557;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_instr <= _GEN_1054;
        end
      end else begin
        REG__6_cf_instr <= _GEN_1054;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_pc <= _GEN_1046;
        end
      end else begin
        REG__6_cf_pc <= _GEN_1046;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_pnpc <= _GEN_1038;
        end
      end else begin
        REG__6_cf_pnpc <= _GEN_1038;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_exceptionVec_1 <= _GEN_894;
        end
      end else begin
        REG__6_cf_exceptionVec_1 <= _GEN_894;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_exceptionVec_2 <= _GEN_902;
        end
      end else begin
        REG__6_cf_exceptionVec_2 <= _GEN_902;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_exceptionVec_12 <= _GEN_982;
        end
      end else begin
        REG__6_cf_exceptionVec_12 <= _GEN_982;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_0 <= _GEN_790;
        end
      end else begin
        REG__6_cf_intrVec_0 <= _GEN_790;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_1 <= _GEN_798;
        end
      end else begin
        REG__6_cf_intrVec_1 <= _GEN_798;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_2 <= _GEN_806;
        end
      end else begin
        REG__6_cf_intrVec_2 <= _GEN_806;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_3 <= _GEN_814;
        end
      end else begin
        REG__6_cf_intrVec_3 <= _GEN_814;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_4 <= _GEN_822;
        end
      end else begin
        REG__6_cf_intrVec_4 <= _GEN_822;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_5 <= _GEN_830;
        end
      end else begin
        REG__6_cf_intrVec_5 <= _GEN_830;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_6 <= _GEN_838;
        end
      end else begin
        REG__6_cf_intrVec_6 <= _GEN_838;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_7 <= _GEN_846;
        end
      end else begin
        REG__6_cf_intrVec_7 <= _GEN_846;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_8 <= _GEN_854;
        end
      end else begin
        REG__6_cf_intrVec_8 <= _GEN_854;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_9 <= _GEN_862;
        end
      end else begin
        REG__6_cf_intrVec_9 <= _GEN_862;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_10 <= _GEN_870;
        end
      end else begin
        REG__6_cf_intrVec_10 <= _GEN_870;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_intrVec_11 <= _GEN_878;
        end
      end else begin
        REG__6_cf_intrVec_11 <= _GEN_878;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_brIdx <= _GEN_782;
        end
      end else begin
        REG__6_cf_brIdx <= _GEN_782;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_crossPageIPFFix <= _GEN_766;
        end
      end else begin
        REG__6_cf_crossPageIPFFix <= _GEN_766;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_runahead_checkpoint_id <= _GEN_758;
        end
      end else begin
        REG__6_cf_runahead_checkpoint_id <= _GEN_758;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_cf_instrType <= _GEN_742;
        end
      end else begin
        REG__6_cf_instrType <= _GEN_742;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__6_ctrl_src1Type <= 3'h6 == _T_20 | _GEN_734;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__6_ctrl_src1Type <= _GEN_206;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__6_ctrl_src2Type <= 3'h6 == _T_20 | _GEN_726;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__6_ctrl_src2Type <= _GEN_198;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_fuType <= _GEN_718;
        end
      end else begin
        REG__6_ctrl_fuType <= _GEN_718;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_fuOpType <= _GEN_710;
        end
      end else begin
        REG__6_ctrl_fuOpType <= _GEN_710;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_funct3 <= _GEN_702;
        end
      end else begin
        REG__6_ctrl_funct3 <= _GEN_702;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_func24 <= _GEN_694;
        end
      end else begin
        REG__6_ctrl_func24 <= _GEN_694;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_func23 <= _GEN_686;
        end
      end else begin
        REG__6_ctrl_func23 <= _GEN_686;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_rfSrc1 <= _GEN_678;
        end
      end else begin
        REG__6_ctrl_rfSrc1 <= _GEN_678;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_rfSrc2 <= _GEN_670;
        end
      end else begin
        REG__6_ctrl_rfSrc2 <= _GEN_670;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_rfSrc3 <= _GEN_662;
        end
      end else begin
        REG__6_ctrl_rfSrc3 <= _GEN_662;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_rfWen <= _GEN_654;
        end
      end else begin
        REG__6_ctrl_rfWen <= _GEN_654;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_rfDest <= _GEN_646;
        end
      end else begin
        REG__6_ctrl_rfDest <= _GEN_646;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_ctrl_isMou <= _GEN_590;
        end
      end else begin
        REG__6_ctrl_isMou <= _GEN_590;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__6_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h6 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__6_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__6_data_imm <= _GEN_558;
        end
      end else begin
        REG__6_data_imm <= _GEN_558;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_instr <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_instr <= _GEN_1055;
        end
      end else begin
        REG__7_cf_instr <= _GEN_1055;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_pc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_pc <= _GEN_1047;
        end
      end else begin
        REG__7_cf_pc <= _GEN_1047;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_pnpc <= 39'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_pnpc <= _GEN_1039;
        end
      end else begin
        REG__7_cf_pnpc <= _GEN_1039;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_exceptionVec_1 <= _GEN_895;
        end
      end else begin
        REG__7_cf_exceptionVec_1 <= _GEN_895;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_exceptionVec_2 <= _GEN_903;
        end
      end else begin
        REG__7_cf_exceptionVec_2 <= _GEN_903;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_exceptionVec_12 <= _GEN_983;
        end
      end else begin
        REG__7_cf_exceptionVec_12 <= _GEN_983;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_0 <= _GEN_791;
        end
      end else begin
        REG__7_cf_intrVec_0 <= _GEN_791;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_1 <= _GEN_799;
        end
      end else begin
        REG__7_cf_intrVec_1 <= _GEN_799;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_2 <= _GEN_807;
        end
      end else begin
        REG__7_cf_intrVec_2 <= _GEN_807;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_3 <= _GEN_815;
        end
      end else begin
        REG__7_cf_intrVec_3 <= _GEN_815;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_4 <= _GEN_823;
        end
      end else begin
        REG__7_cf_intrVec_4 <= _GEN_823;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_5 <= _GEN_831;
        end
      end else begin
        REG__7_cf_intrVec_5 <= _GEN_831;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_6 <= _GEN_839;
        end
      end else begin
        REG__7_cf_intrVec_6 <= _GEN_839;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_7 <= _GEN_847;
        end
      end else begin
        REG__7_cf_intrVec_7 <= _GEN_847;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_8 <= _GEN_855;
        end
      end else begin
        REG__7_cf_intrVec_8 <= _GEN_855;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_9 <= _GEN_863;
        end
      end else begin
        REG__7_cf_intrVec_9 <= _GEN_863;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_10 <= _GEN_871;
        end
      end else begin
        REG__7_cf_intrVec_10 <= _GEN_871;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_intrVec_11 <= _GEN_879;
        end
      end else begin
        REG__7_cf_intrVec_11 <= _GEN_879;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_brIdx <= 4'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_brIdx <= _GEN_783;
        end
      end else begin
        REG__7_cf_brIdx <= _GEN_783;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_crossPageIPFFix <= _GEN_767;
        end
      end else begin
        REG__7_cf_crossPageIPFFix <= _GEN_767;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_runahead_checkpoint_id <= _GEN_759;
        end
      end else begin
        REG__7_cf_runahead_checkpoint_id <= _GEN_759;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_cf_instrType <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_cf_instrType <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_cf_instrType <= _GEN_743;
        end
      end else begin
        REG__7_cf_instrType <= _GEN_743;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__7_ctrl_src1Type <= 3'h7 == _T_20 | _GEN_735;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__7_ctrl_src1Type <= _GEN_207;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        REG__7_ctrl_src2Type <= 3'h7 == _T_20 | _GEN_727;
      end else if (_T_11) begin // @[PipelineVector.scala 45:29]
        REG__7_ctrl_src2Type <= _GEN_199;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_fuType <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_fuType <= 4'h1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_fuType <= _GEN_719;
        end
      end else begin
        REG__7_ctrl_fuType <= _GEN_719;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_fuOpType <= _GEN_711;
        end
      end else begin
        REG__7_ctrl_fuOpType <= _GEN_711;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_funct3 <= 3'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_funct3 <= _GEN_703;
        end
      end else begin
        REG__7_ctrl_funct3 <= _GEN_703;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_func24 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_func24 <= _GEN_695;
        end
      end else begin
        REG__7_ctrl_func24 <= _GEN_695;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_func23 <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_func23 <= _GEN_687;
        end
      end else begin
        REG__7_ctrl_func23 <= _GEN_687;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_rfSrc1 <= _GEN_679;
        end
      end else begin
        REG__7_ctrl_rfSrc1 <= _GEN_679;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_rfSrc2 <= _GEN_671;
        end
      end else begin
        REG__7_ctrl_rfSrc2 <= _GEN_671;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_rfSrc3 <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_rfSrc3 <= _GEN_663;
        end
      end else begin
        REG__7_ctrl_rfSrc3 <= _GEN_663;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_rfWen <= _GEN_655;
        end
      end else begin
        REG__7_ctrl_rfWen <= _GEN_655;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_rfDest <= _GEN_647;
        end
      end else begin
        REG__7_ctrl_rfDest <= _GEN_647;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_ctrl_isMou <= 1'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_ctrl_isMou <= _GEN_591;
        end
      end else begin
        REG__7_ctrl_isMou <= _GEN_591;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__7_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (3'h7 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__7_data_imm <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__7_data_imm <= _GEN_559;
        end
      end else begin
        REG__7_data_imm <= _GEN_559;
      end
    end
    if (reset) begin // @[PipelineVector.scala 30:33]
      REG_1 <= 3'h0; // @[PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[PipelineVector.scala 71:16]
      REG_1 <= 3'h0; // @[PipelineVector.scala 72:24]
    end else if (_T_13) begin // @[PipelineVector.scala 44:14]
      REG_1 <= _T_22; // @[PipelineVector.scala 47:24]
    end
    if (reset) begin // @[PipelineVector.scala 31:33]
      REG_2 <= 3'h0; // @[PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[PipelineVector.scala 71:16]
      REG_2 <= 3'h0; // @[PipelineVector.scala 73:24]
    end else if (_T_35) begin // @[PipelineVector.scala 66:22]
      REG_2 <= _T_37; // @[PipelineVector.scala 67:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG__0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  REG__0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  REG__0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG__0_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG__0_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG__0_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG__0_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG__0_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG__0_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG__0_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG__0_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG__0_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  REG__0_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG__0_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG__0_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG__0_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  REG__0_cf_crossPageIPFFix = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  REG__0_cf_runahead_checkpoint_id = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  REG__0_cf_instrType = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  REG__0_ctrl_src1Type = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  REG__0_ctrl_src2Type = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG__0_ctrl_fuType = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  REG__0_ctrl_fuOpType = _RAND_25[6:0];
  _RAND_26 = {1{`RANDOM}};
  REG__0_ctrl_funct3 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  REG__0_ctrl_func24 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  REG__0_ctrl_func23 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc1 = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc2 = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc3 = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  REG__0_ctrl_rfWen = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  REG__0_ctrl_rfDest = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  REG__0_ctrl_isMou = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  REG__0_data_imm = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  REG__1_cf_instr = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  REG__1_cf_pc = _RAND_37[38:0];
  _RAND_38 = {2{`RANDOM}};
  REG__1_cf_pnpc = _RAND_38[38:0];
  _RAND_39 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_2 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_12 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG__1_cf_intrVec_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG__1_cf_intrVec_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG__1_cf_intrVec_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG__1_cf_intrVec_3 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG__1_cf_intrVec_4 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG__1_cf_intrVec_5 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG__1_cf_intrVec_6 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG__1_cf_intrVec_7 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG__1_cf_intrVec_8 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG__1_cf_intrVec_9 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG__1_cf_intrVec_10 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  REG__1_cf_intrVec_11 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  REG__1_cf_brIdx = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  REG__1_cf_crossPageIPFFix = _RAND_55[0:0];
  _RAND_56 = {2{`RANDOM}};
  REG__1_cf_runahead_checkpoint_id = _RAND_56[63:0];
  _RAND_57 = {1{`RANDOM}};
  REG__1_cf_instrType = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  REG__1_ctrl_src1Type = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  REG__1_ctrl_src2Type = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  REG__1_ctrl_fuType = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  REG__1_ctrl_fuOpType = _RAND_61[6:0];
  _RAND_62 = {1{`RANDOM}};
  REG__1_ctrl_funct3 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  REG__1_ctrl_func24 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  REG__1_ctrl_func23 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc1 = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc2 = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc3 = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  REG__1_ctrl_rfWen = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  REG__1_ctrl_rfDest = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  REG__1_ctrl_isMou = _RAND_70[0:0];
  _RAND_71 = {2{`RANDOM}};
  REG__1_data_imm = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  REG__2_cf_instr = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  REG__2_cf_pc = _RAND_73[38:0];
  _RAND_74 = {2{`RANDOM}};
  REG__2_cf_pnpc = _RAND_74[38:0];
  _RAND_75 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_12 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  REG__2_cf_intrVec_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  REG__2_cf_intrVec_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  REG__2_cf_intrVec_2 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  REG__2_cf_intrVec_3 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  REG__2_cf_intrVec_4 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  REG__2_cf_intrVec_5 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  REG__2_cf_intrVec_6 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  REG__2_cf_intrVec_7 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  REG__2_cf_intrVec_8 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  REG__2_cf_intrVec_9 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  REG__2_cf_intrVec_10 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  REG__2_cf_intrVec_11 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG__2_cf_brIdx = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  REG__2_cf_crossPageIPFFix = _RAND_91[0:0];
  _RAND_92 = {2{`RANDOM}};
  REG__2_cf_runahead_checkpoint_id = _RAND_92[63:0];
  _RAND_93 = {1{`RANDOM}};
  REG__2_cf_instrType = _RAND_93[4:0];
  _RAND_94 = {1{`RANDOM}};
  REG__2_ctrl_src1Type = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  REG__2_ctrl_src2Type = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  REG__2_ctrl_fuType = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  REG__2_ctrl_fuOpType = _RAND_97[6:0];
  _RAND_98 = {1{`RANDOM}};
  REG__2_ctrl_funct3 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  REG__2_ctrl_func24 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG__2_ctrl_func23 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc1 = _RAND_101[4:0];
  _RAND_102 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc2 = _RAND_102[4:0];
  _RAND_103 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc3 = _RAND_103[4:0];
  _RAND_104 = {1{`RANDOM}};
  REG__2_ctrl_rfWen = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  REG__2_ctrl_rfDest = _RAND_105[4:0];
  _RAND_106 = {1{`RANDOM}};
  REG__2_ctrl_isMou = _RAND_106[0:0];
  _RAND_107 = {2{`RANDOM}};
  REG__2_data_imm = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  REG__3_cf_instr = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  REG__3_cf_pc = _RAND_109[38:0];
  _RAND_110 = {2{`RANDOM}};
  REG__3_cf_pnpc = _RAND_110[38:0];
  _RAND_111 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_2 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_12 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG__3_cf_intrVec_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  REG__3_cf_intrVec_1 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  REG__3_cf_intrVec_2 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG__3_cf_intrVec_3 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG__3_cf_intrVec_4 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  REG__3_cf_intrVec_5 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG__3_cf_intrVec_6 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  REG__3_cf_intrVec_7 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  REG__3_cf_intrVec_8 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  REG__3_cf_intrVec_9 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  REG__3_cf_intrVec_10 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  REG__3_cf_intrVec_11 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  REG__3_cf_brIdx = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  REG__3_cf_crossPageIPFFix = _RAND_127[0:0];
  _RAND_128 = {2{`RANDOM}};
  REG__3_cf_runahead_checkpoint_id = _RAND_128[63:0];
  _RAND_129 = {1{`RANDOM}};
  REG__3_cf_instrType = _RAND_129[4:0];
  _RAND_130 = {1{`RANDOM}};
  REG__3_ctrl_src1Type = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  REG__3_ctrl_src2Type = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  REG__3_ctrl_fuType = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  REG__3_ctrl_fuOpType = _RAND_133[6:0];
  _RAND_134 = {1{`RANDOM}};
  REG__3_ctrl_funct3 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  REG__3_ctrl_func24 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  REG__3_ctrl_func23 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc1 = _RAND_137[4:0];
  _RAND_138 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc2 = _RAND_138[4:0];
  _RAND_139 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc3 = _RAND_139[4:0];
  _RAND_140 = {1{`RANDOM}};
  REG__3_ctrl_rfWen = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  REG__3_ctrl_rfDest = _RAND_141[4:0];
  _RAND_142 = {1{`RANDOM}};
  REG__3_ctrl_isMou = _RAND_142[0:0];
  _RAND_143 = {2{`RANDOM}};
  REG__3_data_imm = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  REG__4_cf_instr = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  REG__4_cf_pc = _RAND_145[38:0];
  _RAND_146 = {2{`RANDOM}};
  REG__4_cf_pnpc = _RAND_146[38:0];
  _RAND_147 = {1{`RANDOM}};
  REG__4_cf_exceptionVec_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  REG__4_cf_exceptionVec_2 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  REG__4_cf_exceptionVec_12 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  REG__4_cf_intrVec_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  REG__4_cf_intrVec_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  REG__4_cf_intrVec_2 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  REG__4_cf_intrVec_3 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  REG__4_cf_intrVec_4 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  REG__4_cf_intrVec_5 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  REG__4_cf_intrVec_6 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  REG__4_cf_intrVec_7 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  REG__4_cf_intrVec_8 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  REG__4_cf_intrVec_9 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  REG__4_cf_intrVec_10 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  REG__4_cf_intrVec_11 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  REG__4_cf_brIdx = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  REG__4_cf_crossPageIPFFix = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  REG__4_cf_runahead_checkpoint_id = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  REG__4_cf_instrType = _RAND_165[4:0];
  _RAND_166 = {1{`RANDOM}};
  REG__4_ctrl_src1Type = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  REG__4_ctrl_src2Type = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  REG__4_ctrl_fuType = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  REG__4_ctrl_fuOpType = _RAND_169[6:0];
  _RAND_170 = {1{`RANDOM}};
  REG__4_ctrl_funct3 = _RAND_170[2:0];
  _RAND_171 = {1{`RANDOM}};
  REG__4_ctrl_func24 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  REG__4_ctrl_func23 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  REG__4_ctrl_rfSrc1 = _RAND_173[4:0];
  _RAND_174 = {1{`RANDOM}};
  REG__4_ctrl_rfSrc2 = _RAND_174[4:0];
  _RAND_175 = {1{`RANDOM}};
  REG__4_ctrl_rfSrc3 = _RAND_175[4:0];
  _RAND_176 = {1{`RANDOM}};
  REG__4_ctrl_rfWen = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  REG__4_ctrl_rfDest = _RAND_177[4:0];
  _RAND_178 = {1{`RANDOM}};
  REG__4_ctrl_isMou = _RAND_178[0:0];
  _RAND_179 = {2{`RANDOM}};
  REG__4_data_imm = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  REG__5_cf_instr = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  REG__5_cf_pc = _RAND_181[38:0];
  _RAND_182 = {2{`RANDOM}};
  REG__5_cf_pnpc = _RAND_182[38:0];
  _RAND_183 = {1{`RANDOM}};
  REG__5_cf_exceptionVec_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  REG__5_cf_exceptionVec_2 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  REG__5_cf_exceptionVec_12 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  REG__5_cf_intrVec_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  REG__5_cf_intrVec_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  REG__5_cf_intrVec_2 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  REG__5_cf_intrVec_3 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  REG__5_cf_intrVec_4 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  REG__5_cf_intrVec_5 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  REG__5_cf_intrVec_6 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  REG__5_cf_intrVec_7 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  REG__5_cf_intrVec_8 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  REG__5_cf_intrVec_9 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  REG__5_cf_intrVec_10 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  REG__5_cf_intrVec_11 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  REG__5_cf_brIdx = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  REG__5_cf_crossPageIPFFix = _RAND_199[0:0];
  _RAND_200 = {2{`RANDOM}};
  REG__5_cf_runahead_checkpoint_id = _RAND_200[63:0];
  _RAND_201 = {1{`RANDOM}};
  REG__5_cf_instrType = _RAND_201[4:0];
  _RAND_202 = {1{`RANDOM}};
  REG__5_ctrl_src1Type = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  REG__5_ctrl_src2Type = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  REG__5_ctrl_fuType = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  REG__5_ctrl_fuOpType = _RAND_205[6:0];
  _RAND_206 = {1{`RANDOM}};
  REG__5_ctrl_funct3 = _RAND_206[2:0];
  _RAND_207 = {1{`RANDOM}};
  REG__5_ctrl_func24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  REG__5_ctrl_func23 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  REG__5_ctrl_rfSrc1 = _RAND_209[4:0];
  _RAND_210 = {1{`RANDOM}};
  REG__5_ctrl_rfSrc2 = _RAND_210[4:0];
  _RAND_211 = {1{`RANDOM}};
  REG__5_ctrl_rfSrc3 = _RAND_211[4:0];
  _RAND_212 = {1{`RANDOM}};
  REG__5_ctrl_rfWen = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  REG__5_ctrl_rfDest = _RAND_213[4:0];
  _RAND_214 = {1{`RANDOM}};
  REG__5_ctrl_isMou = _RAND_214[0:0];
  _RAND_215 = {2{`RANDOM}};
  REG__5_data_imm = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  REG__6_cf_instr = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  REG__6_cf_pc = _RAND_217[38:0];
  _RAND_218 = {2{`RANDOM}};
  REG__6_cf_pnpc = _RAND_218[38:0];
  _RAND_219 = {1{`RANDOM}};
  REG__6_cf_exceptionVec_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  REG__6_cf_exceptionVec_2 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  REG__6_cf_exceptionVec_12 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  REG__6_cf_intrVec_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  REG__6_cf_intrVec_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  REG__6_cf_intrVec_2 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  REG__6_cf_intrVec_3 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  REG__6_cf_intrVec_4 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  REG__6_cf_intrVec_5 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  REG__6_cf_intrVec_6 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  REG__6_cf_intrVec_7 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  REG__6_cf_intrVec_8 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  REG__6_cf_intrVec_9 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  REG__6_cf_intrVec_10 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  REG__6_cf_intrVec_11 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  REG__6_cf_brIdx = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  REG__6_cf_crossPageIPFFix = _RAND_235[0:0];
  _RAND_236 = {2{`RANDOM}};
  REG__6_cf_runahead_checkpoint_id = _RAND_236[63:0];
  _RAND_237 = {1{`RANDOM}};
  REG__6_cf_instrType = _RAND_237[4:0];
  _RAND_238 = {1{`RANDOM}};
  REG__6_ctrl_src1Type = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  REG__6_ctrl_src2Type = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  REG__6_ctrl_fuType = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  REG__6_ctrl_fuOpType = _RAND_241[6:0];
  _RAND_242 = {1{`RANDOM}};
  REG__6_ctrl_funct3 = _RAND_242[2:0];
  _RAND_243 = {1{`RANDOM}};
  REG__6_ctrl_func24 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  REG__6_ctrl_func23 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  REG__6_ctrl_rfSrc1 = _RAND_245[4:0];
  _RAND_246 = {1{`RANDOM}};
  REG__6_ctrl_rfSrc2 = _RAND_246[4:0];
  _RAND_247 = {1{`RANDOM}};
  REG__6_ctrl_rfSrc3 = _RAND_247[4:0];
  _RAND_248 = {1{`RANDOM}};
  REG__6_ctrl_rfWen = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  REG__6_ctrl_rfDest = _RAND_249[4:0];
  _RAND_250 = {1{`RANDOM}};
  REG__6_ctrl_isMou = _RAND_250[0:0];
  _RAND_251 = {2{`RANDOM}};
  REG__6_data_imm = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  REG__7_cf_instr = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  REG__7_cf_pc = _RAND_253[38:0];
  _RAND_254 = {2{`RANDOM}};
  REG__7_cf_pnpc = _RAND_254[38:0];
  _RAND_255 = {1{`RANDOM}};
  REG__7_cf_exceptionVec_1 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  REG__7_cf_exceptionVec_2 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  REG__7_cf_exceptionVec_12 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  REG__7_cf_intrVec_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  REG__7_cf_intrVec_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  REG__7_cf_intrVec_2 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  REG__7_cf_intrVec_3 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  REG__7_cf_intrVec_4 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  REG__7_cf_intrVec_5 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  REG__7_cf_intrVec_6 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  REG__7_cf_intrVec_7 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  REG__7_cf_intrVec_8 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  REG__7_cf_intrVec_9 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  REG__7_cf_intrVec_10 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  REG__7_cf_intrVec_11 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  REG__7_cf_brIdx = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  REG__7_cf_crossPageIPFFix = _RAND_271[0:0];
  _RAND_272 = {2{`RANDOM}};
  REG__7_cf_runahead_checkpoint_id = _RAND_272[63:0];
  _RAND_273 = {1{`RANDOM}};
  REG__7_cf_instrType = _RAND_273[4:0];
  _RAND_274 = {1{`RANDOM}};
  REG__7_ctrl_src1Type = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  REG__7_ctrl_src2Type = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  REG__7_ctrl_fuType = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  REG__7_ctrl_fuOpType = _RAND_277[6:0];
  _RAND_278 = {1{`RANDOM}};
  REG__7_ctrl_funct3 = _RAND_278[2:0];
  _RAND_279 = {1{`RANDOM}};
  REG__7_ctrl_func24 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  REG__7_ctrl_func23 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  REG__7_ctrl_rfSrc1 = _RAND_281[4:0];
  _RAND_282 = {1{`RANDOM}};
  REG__7_ctrl_rfSrc2 = _RAND_282[4:0];
  _RAND_283 = {1{`RANDOM}};
  REG__7_ctrl_rfSrc3 = _RAND_283[4:0];
  _RAND_284 = {1{`RANDOM}};
  REG__7_ctrl_rfWen = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  REG__7_ctrl_rfDest = _RAND_285[4:0];
  _RAND_286 = {1{`RANDOM}};
  REG__7_ctrl_isMou = _RAND_286[0:0];
  _RAND_287 = {2{`RANDOM}};
  REG__7_data_imm = _RAND_287[63:0];
  _RAND_288 = {1{`RANDOM}};
  REG_1 = _RAND_288[2:0];
  _RAND_289 = {1{`RANDOM}};
  REG_2 = _RAND_289[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  output        io_out_mem_resp_ready,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_out_coh_req_ready,
  output        io_out_coh_req_valid,
  output [31:0] io_out_coh_req_bits_addr,
  output [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_ready,
  input         io_out_coh_resp_valid,
  input  [3:0]  io_out_coh_resp_bits_cmd,
  input  [63:0] io_out_coh_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[Coherence.scala 46:24]
  wire  _T_1 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_14 = ~inflight; // @[Coherence.scala 52:42]
  wire  _T_20 = ~inflight & _T_4; // @[Coherence.scala 52:52]
  reg [31:0] reqLatch_addr; // @[Reg.scala 15:16]
  reg [3:0] reqLatch_cmd; // @[Reg.scala 15:16]
  reg [63:0] reqLatch_wdata; // @[Reg.scala 15:16]
  wire  _T_23 = io_in_req_valid & _T_14; // @[Coherence.scala 65:43]
  wire  _GEN_5 = _T_4 & _T_23; // @[Coherence.scala 63:24 67:39 68:26]
  wire  _GEN_6 = _T_4 & (io_out_coh_req_ready & _T_14); // @[Coherence.scala 62:17 67:39 69:19]
  wire  _GEN_7 = io_in_req_bits_cmd[0] & (io_in_req_valid & _T_14); // @[Coherence.scala 61:24 64:61 65:26]
  wire  _T_36 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_43 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [2:0] _GEN_10 = _T_43 ? 3'h5 : state; // @[Coherence.scala 45:22 78:{48,56}]
  wire  _T_45 = io_out_coh_resp_ready & io_out_coh_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_46 = io_out_coh_resp_bits_cmd == 4'hc; // @[SimpleBus.scala 92:26]
  wire [2:0] _T_47 = _T_46 ? 3'h2 : 3'h3; // @[Coherence.scala 83:21]
  wire  _T_50 = io_in_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [2:0] _GEN_14 = io_in_resp_valid & _T_50 ? 3'h0 : state; // @[Coherence.scala 45:22 89:{60,68}]
  wire  _T_53 = io_out_mem_req_ready & io_out_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_53 ? 3'h4 : state; // @[Coherence.scala 45:22 94:{36,44}]
  wire  _T_55 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_56 = io_out_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [2:0] _GEN_16 = _T_55 & _T_56 ? 3'h0 : state; // @[Coherence.scala 96:101 45:22 96:93]
  wire [2:0] _GEN_17 = _T_55 ? 3'h0 : state; // @[Coherence.scala 45:22 97:{57,65}]
  wire [2:0] _GEN_18 = 3'h5 == state ? _GEN_17 : state; // @[Coherence.scala 74:18 45:22]
  wire [2:0] _GEN_19 = 3'h4 == state ? _GEN_16 : _GEN_18; // @[Coherence.scala 74:18]
  wire [63:0] _GEN_20 = 3'h3 == state ? reqLatch_wdata : io_in_req_bits_wdata; // @[Coherence.scala 74:18 59:23 92:27]
  wire [3:0] _GEN_22 = 3'h3 == state ? reqLatch_cmd : io_in_req_bits_cmd; // @[Coherence.scala 74:18 59:23 92:27]
  wire [31:0] _GEN_24 = 3'h3 == state ? reqLatch_addr : io_in_req_bits_addr; // @[Coherence.scala 74:18 59:23 92:27]
  wire  _GEN_25 = 3'h3 == state | _GEN_7; // @[Coherence.scala 74:18 93:28]
  wire [2:0] _GEN_26 = 3'h3 == state ? _GEN_15 : _GEN_19; // @[Coherence.scala 74:18]
  wire [63:0] _GEN_27 = 3'h2 == state ? io_out_coh_resp_bits_rdata : io_out_mem_resp_bits_rdata; // @[Coherence.scala 72:14 74:18 88:16]
  wire [3:0] _GEN_28 = 3'h2 == state ? io_out_coh_resp_bits_cmd : io_out_mem_resp_bits_cmd; // @[Coherence.scala 72:14 74:18 88:16]
  wire  _GEN_29 = 3'h2 == state ? io_out_coh_resp_valid : io_out_mem_resp_valid; // @[Coherence.scala 72:14 74:18 88:16]
  wire [63:0] _GEN_32 = 3'h2 == state ? io_in_req_bits_wdata : _GEN_20; // @[Coherence.scala 74:18 59:23]
  wire [3:0] _GEN_34 = 3'h2 == state ? io_in_req_bits_cmd : _GEN_22; // @[Coherence.scala 74:18 59:23]
  wire [31:0] _GEN_36 = 3'h2 == state ? io_in_req_bits_addr : _GEN_24; // @[Coherence.scala 74:18 59:23]
  wire  _GEN_37 = 3'h2 == state ? _GEN_7 : _GEN_25; // @[Coherence.scala 74:18]
  wire [63:0] _GEN_39 = 3'h1 == state ? io_out_mem_resp_bits_rdata : _GEN_27; // @[Coherence.scala 72:14 74:18]
  wire [3:0] _GEN_40 = 3'h1 == state ? io_out_mem_resp_bits_cmd : _GEN_28; // @[Coherence.scala 72:14 74:18]
  wire  _GEN_41 = 3'h1 == state ? io_out_mem_resp_valid : _GEN_29; // @[Coherence.scala 72:14 74:18]
  wire [63:0] _GEN_43 = 3'h1 == state ? io_in_req_bits_wdata : _GEN_32; // @[Coherence.scala 74:18 59:23]
  wire [3:0] _GEN_45 = 3'h1 == state ? io_in_req_bits_cmd : _GEN_34; // @[Coherence.scala 74:18 59:23]
  wire [31:0] _GEN_47 = 3'h1 == state ? io_in_req_bits_addr : _GEN_36; // @[Coherence.scala 74:18 59:23]
  wire  _GEN_48 = 3'h1 == state ? _GEN_7 : _GEN_37; // @[Coherence.scala 74:18]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? io_out_mem_req_ready & _T_14 : _GEN_6; // @[Coherence.scala 64:61 66:19]
  assign io_in_resp_valid = 3'h0 == state ? io_out_mem_resp_valid : _GEN_41; // @[Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_cmd = 3'h0 == state ? io_out_mem_resp_bits_cmd : _GEN_40; // @[Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_rdata = 3'h0 == state ? io_out_mem_resp_bits_rdata : _GEN_39; // @[Coherence.scala 72:14 74:18]
  assign io_out_mem_req_valid = 3'h0 == state ? _GEN_7 : _GEN_48; // @[Coherence.scala 74:18]
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_47; // @[Coherence.scala 74:18 59:23]
  assign io_out_mem_req_bits_cmd = 3'h0 == state ? io_in_req_bits_cmd : _GEN_45; // @[Coherence.scala 74:18 59:23]
  assign io_out_mem_req_bits_wdata = 3'h0 == state ? io_in_req_bits_wdata : _GEN_43; // @[Coherence.scala 74:18 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[Coherence.scala 72:14]
  assign io_out_coh_req_valid = io_in_req_bits_cmd[0] ? 1'h0 : _GEN_5; // @[Coherence.scala 63:24 64:61]
  assign io_out_coh_req_bits_addr = io_in_req_bits_addr; // @[Coherence.scala 54:16]
  assign io_out_coh_req_bits_wdata = io_in_req_bits_wdata; // @[Coherence.scala 54:16]
  assign io_out_coh_resp_ready = 1'h1; // @[Coherence.scala 56:18 74:18]
  always @(posedge clock) begin
    if (reset) begin // @[Coherence.scala 45:22]
      state <= 3'h0; // @[Coherence.scala 45:22]
    end else if (3'h0 == state) begin // @[Coherence.scala 74:18]
      if (_T_36) begin // @[Coherence.scala 76:29]
        if (_T_4) begin // @[Coherence.scala 77:38]
          state <= 3'h1; // @[Coherence.scala 77:46]
        end else begin
          state <= _GEN_10;
        end
      end
    end else if (3'h1 == state) begin // @[Coherence.scala 74:18]
      if (_T_45) begin // @[Coherence.scala 82:37]
        state <= _T_47; // @[Coherence.scala 83:15]
      end
    end else if (3'h2 == state) begin // @[Coherence.scala 74:18]
      state <= _GEN_14;
    end else begin
      state <= _GEN_26;
    end
    if (_T_20) begin // @[Reg.scala 16:19]
      reqLatch_addr <= io_in_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (_T_20) begin // @[Reg.scala 16:19]
      reqLatch_cmd <= io_in_req_bits_cmd; // @[Reg.scala 16:23]
    end
    if (_T_20) begin // @[Reg.scala 16:19]
      reqLatch_wdata <= io_in_req_bits_wdata; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Coherence.scala:49 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Coherence.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Coherence.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_cmd = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  reqLatch_wdata = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI42SimpleBusConverter(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  input  [17:0] io_in_awid,
  input  [7:0]  io_in_awlen,
  input  [2:0]  io_in_awsize,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_wlast,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input  [17:0] io_in_arid,
  input  [7:0]  io_in_arlen,
  input  [2:0]  io_in_arsize,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata,
  output        io_in_rlast,
  output [17:0] io_in_rid,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] inflight_id_reg; // @[ToAXI4.scala 38:32]
  reg [1:0] inflight_type; // @[ToAXI4.scala 40:30]
  wire  _T = inflight_type == 2'h0; // @[ToAXI4.scala 50:19]
  wire  _T_1 = ~_T; // @[ToAXI4.scala 53:5]
  wire  _T_2 = ~_T_1; // @[ToAXI4.scala 64:9]
  wire  _T_3 = ~_T_1 & io_in_arvalid; // @[ToAXI4.scala 64:23]
  wire [1:0] _T_5 = io_in_arlen == 8'h0 ? 2'h0 : 2'h2; // @[ToAXI4.scala 67:19]
  wire  _T_6 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [17:0] _GEN_0 = _T_6 ? io_in_arid : inflight_id_reg; // @[ToAXI4.scala 42:21 74:25 38:32]
  wire [1:0] _GEN_1 = _T_6 ? 2'h1 : inflight_type; // @[ToAXI4.scala 43:19 74:25 40:30]
  wire [31:0] _GEN_2 = ~_T_1 & io_in_arvalid ? io_in_araddr : 32'h0; // @[ToAXI4.scala 64:40 66:14 59:7]
  wire [3:0] _GEN_3 = ~_T_1 & io_in_arvalid ? {{2'd0}, _T_5} : 4'h0; // @[ToAXI4.scala 64:40 67:13 59:7]
  wire [2:0] _GEN_4 = ~_T_1 & io_in_arvalid ? io_in_arsize : 3'h0; // @[ToAXI4.scala 64:40 69:14 59:7]
  wire [17:0] _GEN_7 = ~_T_1 & io_in_arvalid ? _GEN_0 : inflight_id_reg; // @[ToAXI4.scala 38:32 64:40]
  wire [1:0] _GEN_8 = ~_T_1 & io_in_arvalid ? _GEN_1 : inflight_type; // @[ToAXI4.scala 40:30 64:40]
  wire  _T_7 = inflight_type == 2'h1; // @[ToAXI4.scala 50:19]
  wire  _T_9 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_10 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_9 = _T_10 & _T_9 ? 2'h0 : _GEN_8; // @[ToAXI4.scala 46:19 88:42]
  wire [17:0] _GEN_10 = _T_10 & _T_9 ? 18'h0 : _GEN_7; // @[ToAXI4.scala 47:21 88:42]
  wire [1:0] _GEN_15 = _T_7 & io_out_resp_valid ? _GEN_9 : _GEN_8; // @[ToAXI4.scala 79:46]
  wire [17:0] _GEN_16 = _T_7 & io_out_resp_valid ? _GEN_10 : _GEN_7; // @[ToAXI4.scala 79:46]
  reg [31:0] aw_reg_addr; // @[ToAXI4.scala 94:19]
  reg [7:0] aw_reg_len; // @[ToAXI4.scala 94:19]
  reg [2:0] aw_reg_size; // @[ToAXI4.scala 94:19]
  reg  bresp_en; // @[ToAXI4.scala 95:25]
  wire  _T_17 = ~io_in_arvalid; // @[ToAXI4.scala 97:42]
  wire  _T_19 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_20 = inflight_type == 2'h2; // @[ToAXI4.scala 50:19]
  wire  _T_21 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_24 = io_in_wlast ? 3'h7 : 3'h3; // @[ToAXI4.scala 108:10]
  wire [2:0] _T_25 = aw_reg_len == 8'h0 ? 3'h1 : _T_24; // @[ToAXI4.scala 107:19]
  wire  _GEN_31 = io_in_wlast | bresp_en; // @[ToAXI4.scala 115:19 116:16 95:25]
  wire  _T_26 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  wire  _T_57 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_81 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  assign io_in_awready = _T_2 & _T_17; // @[ToAXI4.scala 132:33]
  assign io_in_wready = _T_20 & io_out_req_ready; // @[ToAXI4.scala 133:38]
  assign io_in_bvalid = bresp_en & io_out_resp_valid; // @[ToAXI4.scala 134:27]
  assign io_in_arready = _T_2 & io_out_req_ready; // @[ToAXI4.scala 129:33]
  assign io_in_rvalid = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 130:36]
  assign io_in_rdata = _T_7 & io_out_resp_valid ? io_out_resp_bits_rdata : 64'h0; // @[ToAXI4.scala 79:46 81:12 60:5]
  assign io_in_rlast = _T_7 & io_out_resp_valid & _T_9; // @[ToAXI4.scala 79:46 85:12 60:5]
  assign io_in_rid = _T_7 & io_out_resp_valid ? inflight_id_reg : 18'h0; // @[ToAXI4.scala 79:46 82:10 60:5]
  assign io_out_req_valid = _T_3 | _T_20 & io_in_wvalid; // @[ToAXI4.scala 127:52]
  assign io_out_req_bits_addr = _T_20 & _T_21 ? aw_reg_addr : _GEN_2; // @[ToAXI4.scala 105:45 109:14]
  assign io_out_req_bits_size = _T_20 & _T_21 ? aw_reg_size : _GEN_4; // @[ToAXI4.scala 105:45 110:14]
  assign io_out_req_bits_cmd = _T_20 & _T_21 ? {{1'd0}, _T_25} : _GEN_3; // @[ToAXI4.scala 105:45 107:13]
  assign io_out_req_bits_wmask = _T_20 & _T_21 ? io_in_wstrb : 8'h0; // @[ToAXI4.scala 105:45 111:15]
  assign io_out_req_bits_wdata = _T_20 & _T_21 ? io_in_wdata : 64'h0; // @[ToAXI4.scala 105:45 112:15]
  assign io_out_resp_ready = _T_2 | _T_7 & io_in_rready | _T_20 & io_in_bready; // @[ToAXI4.scala 128:73]
  always @(posedge clock) begin
    if (reset) begin // @[ToAXI4.scala 38:32]
      inflight_id_reg <= 18'h0; // @[ToAXI4.scala 38:32]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      inflight_id_reg <= 18'h0; // @[ToAXI4.scala 47:21]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      if (_T_19) begin // @[ToAXI4.scala 100:24]
        inflight_id_reg <= io_in_awid; // @[ToAXI4.scala 42:21]
      end else begin
        inflight_id_reg <= _GEN_16;
      end
    end else begin
      inflight_id_reg <= _GEN_16;
    end
    if (reset) begin // @[ToAXI4.scala 40:30]
      inflight_type <= 2'h0; // @[ToAXI4.scala 40:30]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      inflight_type <= 2'h0; // @[ToAXI4.scala 46:19]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      if (_T_19) begin // @[ToAXI4.scala 100:24]
        inflight_type <= 2'h2; // @[ToAXI4.scala 43:19]
      end else begin
        inflight_type <= _GEN_15;
      end
    end else begin
      inflight_type <= _GEN_15;
    end
    if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_addr <= io_in_awaddr; // @[ToAXI4.scala 98:12]
    end
    if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_len <= io_in_awlen; // @[ToAXI4.scala 98:12]
    end
    if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_size <= io_in_awsize; // @[ToAXI4.scala 98:12]
    end
    if (reset) begin // @[ToAXI4.scala 95:25]
      bresp_en <= 1'h0; // @[ToAXI4.scala 95:25]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      bresp_en <= 1'h0; // @[ToAXI4.scala 121:14]
    end else if (_T_20 & _T_21) begin // @[ToAXI4.scala 105:45]
      bresp_en <= _GEN_31;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & ~(_T_6 & _T_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:137 when (axi.ar.fire()) { assert(mem.req.fire() && !isInflight()); }\n"
            ); // @[ToAXI4.scala 137:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_57 & ~(_T_6 & _T_2 | reset)) begin
          $fatal; // @[ToAXI4.scala 137:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & ~(_T_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:138 when (axi.aw.fire()) { assert(!isInflight()); }\n"); // @[ToAXI4.scala 138:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_19 & ~(_T_2 | reset)) begin
          $fatal; // @[ToAXI4.scala 138:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & ~(_T_6 & _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:139 when (axi.w.fire()) { assert(mem.req .fire() && isState(axi_write)); }\n"
            ); // @[ToAXI4.scala 139:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21 & ~(_T_6 & _T_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 139:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26 & ~(_T_81 & _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:140 when (axi.b.fire()) { assert(mem.resp.fire() && isState(axi_write)); }\n"
            ); // @[ToAXI4.scala 140:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_26 & ~(_T_81 & _T_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 140:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(_T_81 & _T_7 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:141 when (axi.r.fire()) { assert(mem.resp.fire() && isState(axi_read)); }\n"
            ); // @[ToAXI4.scala 141:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10 & ~(_T_81 & _T_7 | reset)) begin
          $fatal; // @[ToAXI4.scala 141:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inflight_id_reg = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  inflight_type = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  aw_reg_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  aw_reg_len = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  aw_reg_size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bresp_en = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Prefetcher(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  getNewReq; // @[Prefetcher.scala 37:26]
  reg [31:0] prefetchReq_addr; // @[Prefetcher.scala 38:28]
  reg [2:0] prefetchReq_size; // @[Prefetcher.scala 38:28]
  reg [7:0] prefetchReq_wmask; // @[Prefetcher.scala 38:28]
  reg [63:0] prefetchReq_wdata; // @[Prefetcher.scala 38:28]
  reg [63:0] lastReqAddr; // @[Prefetcher.scala 44:28]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_9 = {{32'd0}, io_in_bits_addr}; // @[Prefetcher.scala 50:30]
  wire [63:0] _T_4 = _GEN_9 & 64'hffffffffffffffc0; // @[Prefetcher.scala 50:30]
  wire [63:0] _T_5 = lastReqAddr & 64'hffffffffffffffc0; // @[Prefetcher.scala 50:59]
  wire  neqAddr = _T_4 != _T_5; // @[Prefetcher.scala 50:42]
  wire  _T_8 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = prefetchReq_addr < 32'h40000000; // @[NutCore.scala 92:35]
  wire  _T_19 = prefetchReq_addr >= 32'h40600000 & prefetchReq_addr < 32'h41600000; // @[NutCore.scala 92:26]
  wire  _T_20 = _T_15 | _T_19; // @[NutCore.scala 93:15]
  assign io_in_ready = ~getNewReq & (~io_in_valid | _T_8); // @[Prefetcher.scala 52:21 55:17 60:17]
  assign io_out_valid = ~getNewReq ? io_in_valid : ~_T_20; // @[Prefetcher.scala 52:21 54:18 59:18]
  assign io_out_bits_addr = ~getNewReq ? io_in_bits_addr : prefetchReq_addr; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_size = ~getNewReq ? io_in_bits_size : prefetchReq_size; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_cmd = ~getNewReq ? io_in_bits_cmd : 4'h4; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_wmask = ~getNewReq ? io_in_bits_wmask : prefetchReq_wmask; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_wdata = ~getNewReq ? io_in_bits_wdata : prefetchReq_wdata; // @[Prefetcher.scala 52:21 53:17 58:17]
  always @(posedge clock) begin
    if (reset) begin // @[Prefetcher.scala 37:26]
      getNewReq <= 1'h0; // @[Prefetcher.scala 37:26]
    end else if (~getNewReq) begin // @[Prefetcher.scala 52:21]
      getNewReq <= _T_2 & io_in_bits_cmd[1] & neqAddr; // @[Prefetcher.scala 56:15]
    end else begin
      getNewReq <= ~(_T_8 | _T_20); // @[Prefetcher.scala 61:15]
    end
    prefetchReq_addr <= io_in_bits_addr + 32'h40; // @[Prefetcher.scala 40:39]
    prefetchReq_size <= io_in_bits_size; // @[Prefetcher.scala 38:28]
    prefetchReq_wmask <= io_in_bits_wmask; // @[Prefetcher.scala 38:28]
    prefetchReq_wdata <= io_in_bits_wdata; // @[Prefetcher.scala 38:28]
    if (reset) begin // @[Prefetcher.scala 44:28]
      lastReqAddr <= 64'h0; // @[Prefetcher.scala 44:28]
    end else if (_T_2) begin // @[Prefetcher.scala 45:23]
      lastReqAddr <= {{32'd0}, io_in_bits_addr}; // @[Prefetcher.scala 46:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  getNewReq = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  prefetchReq_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  prefetchReq_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  prefetchReq_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  prefetchReq_wdata = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  lastReqAddr = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1_2(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [8:0]  io_metaReadBus_req_bits_setIdx,
  input  [16:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [16:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [16:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [16:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_24 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_24) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 147:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 146:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 145:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 145:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 145:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 145:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[14:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[14:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module CacheStage2_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [16:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_dirty,
  output [16:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_dirty,
  output [16:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_dirty,
  output [16:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [16:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [16:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [16:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [16:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [8:0]  io_metaWriteBus_req_bits_setIdx,
  input  [16:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [11:0] io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 176:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 176:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 176:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 178:64]
  reg  isForwardMetaReg; // @[Cache.scala 179:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 180:24 179:33 180:43]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 181:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 181:22]
  reg [16:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 15:16 16:{19,23}]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 15:16 16:{19,23}]
  wire [16:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 15:16 16:{19,23}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 185:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 187:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 187:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 187:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 187:61]
  wire [16:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[Cache.scala 189:22]
  wire [16:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[Cache.scala 189:22]
  wire [16:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[Cache.scala 189:22]
  wire [16:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[Cache.scala 189:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 192:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_39 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_42 = {_T_39,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 193:42]
  wire  _T_45 = ~metaWay_0_valid; // @[Cache.scala 195:45]
  wire  _T_46 = ~metaWay_1_valid; // @[Cache.scala 195:45]
  wire  _T_47 = ~metaWay_2_valid; // @[Cache.scala 195:45]
  wire  _T_48 = ~metaWay_3_valid; // @[Cache.scala 195:45]
  wire [3:0] invalidVec = {_T_48,_T_47,_T_46,_T_45}; // @[Cache.scala 195:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 196:34]
  wire [1:0] _T_52 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 199:8]
  wire [2:0] _T_53 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_52}; // @[Cache.scala 198:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_53}; // @[Cache.scala 197:33]
  wire [3:0] _T_54 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 202:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  wire [1:0] _T_59 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_61 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_63 = _T_59 + _T_61; // @[Bitwise.scala 47:55]
  wire  _T_65 = _T_63 > 3'h1; // @[Cache.scala 203:26]
  wire  _T_173 = io_in_bits_req_addr < 32'h40000000; // @[NutCore.scala 92:35]
  wire  _T_177 = io_in_bits_req_addr >= 32'h40600000 & io_in_bits_req_addr < 32'h41600000; // @[NutCore.scala 92:26]
  wire [11:0] _T_194 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_196 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_194; // @[Cache.scala 220:13]
  wire  isForwardData = io_in_valid & _T_196; // @[Cache.scala 219:35]
  reg  isForwardDataReg; // @[Cache.scala 222:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 223:24 222:33 223:43]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_203 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_203; // @[Cache.scala 231:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 230:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 229:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 229:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 229:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 229:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 215:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 213:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  assign io_out_bits_mmio = _T_173 | _T_177; // @[NutCore.scala 93:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 226:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 227:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 227:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 179:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 179:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 181:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 181:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_42;
    end
    if (reset) begin // @[Cache.scala 222:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 222:33]
    end else if (_T_12) begin // @[Cache.scala 224:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 224:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 16:23]
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:210 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 210:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fatal; // @[Cache.scala 210:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  REG = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_10(
  input         io_in_0_valid,
  input  [8:0]  io_in_0_bits_setIdx,
  input  [16:0] io_in_0_bits_data_tag,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [8:0]  io_in_1_bits_setIdx,
  input  [16:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [8:0]  io_out_bits_setIdx,
  output [16:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid | io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module Arbiter_11(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module CacheStage3_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [16:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_dirty,
  input  [16:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_dirty,
  input  [16:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_dirty,
  input  [16:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [11:0] io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [8:0]  io_metaWriteBus_req_bits_setIdx,
  output [16:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  output        io_cohResp_valid,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 257:28]
  wire [8:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 257:28]
  wire [16:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 257:28]
  wire [8:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 257:28]
  wire [16:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 257:28]
  wire [8:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 257:28]
  wire [16:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 257:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 257:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 258:28]
  wire [11:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 258:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 258:28]
  wire [11:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 258:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 258:28]
  wire [11:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 258:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 258:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 258:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 261:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 261:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 262:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 263:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 264:26]
  wire  _T_6 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_6; // @[Cache.scala 265:39]
  wire  _T_7 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_7; // @[Cache.scala 266:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[Mux.scala 27:72]
  wire [16:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [16:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [16:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 277:49]
  wire [63:0] _T_50 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_51 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_52 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_53 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_54 = _T_50 | _T_51; // @[Mux.scala 27:72]
  wire [63:0] _T_55 = _T_54 | _T_52; // @[Mux.scala 27:72]
  wire [63:0] _T_56 = _T_55 | _T_53; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_56; // @[Cache.scala 279:21]
  wire [7:0] _T_69 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_77 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_79 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_81 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_83 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_84 = {_T_83,_T_81,_T_79,_T_77,_T_75,_T_73,_T_71,_T_69}; // @[Cat.scala 30:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_84 : 64'h0; // @[Cache.scala 280:21]
  reg [2:0] value; // @[Counter.scala 60:40]
  wire  _T_86 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 283:34]
  wire  _T_87 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_88 = io_in_bits_req_cmd == 4'h3 | _T_87; // @[Cache.scala 283:62]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_0 = io_out_valid & (io_in_bits_req_cmd == 4'h3 | _T_87) ? _value_T_1 : value; // @[Cache.scala 283:85 Counter.scala 76:15 60:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 287:22]
  wire [63:0] _T_91 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_92 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_93 = dataRead & _T_92; // @[BitUtils.scala 32:36]
  wire [2:0] _T_98 = _T_88 ? value : addr_wordIndex; // @[Cache.scala 290:51]
  wire  metaHitWriteBus_req_valid = hitWrite & ~meta_dirty; // @[Cache.scala 293:22]
  reg [3:0] state; // @[Cache.scala 298:22]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 308:23]
  wire  _T_110 = state == 4'h3; // @[Cache.scala 310:39]
  wire  _T_111 = state == 4'h8; // @[Cache.scala 310:66]
  wire [2:0] _T_116 = _T_111 ? value_1 : value_2; // @[Cache.scala 311:33]
  wire  _T_118 = state2 == 2'h1; // @[Cache.scala 312:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_123 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_124 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_125 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_126 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_127 = _T_123 | _T_124; // @[Mux.scala 27:72]
  wire [63:0] _T_128 = _T_127 | _T_125; // @[Mux.scala 27:72]
  wire [63:0] _T_129 = _T_128 | _T_126; // @[Mux.scala 27:72]
  wire  _T_131 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_134 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_8 = _T_134 | io_cohResp_valid | hitReadBurst ? 2'h0 : state2; // @[Cache.scala 318:{100,109} 308:23]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_140 = state == 4'h1; // @[Cache.scala 326:23]
  wire [2:0] _T_142 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 327:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_142; // @[Cache.scala 326:16]
  wire  _T_148 = state2 == 2'h2; // @[Cache.scala 333:89]
  reg  afterFirstRead; // @[Cache.scala 340:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = io_out_valid | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_154 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_156 = state == 4'h2; // @[Cache.scala 342:70]
  wire  readingFirst = ~afterFirstRead & _T_154 & state == 4'h2; // @[Cache.scala 342:60]
  wire  _T_159 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 344:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_160 = state == 4'h0; // @[Cache.scala 347:31]
  wire  _T_164 = _T_111 & _T_148; // @[Cache.scala 348:46]
  wire  _T_168 = _T_111 & io_cohResp_valid; // @[Cache.scala 350:49]
  reg [2:0] value_3; // @[Counter.scala 60:40]
  wire  wrap_wrap = value_3 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_1 = value_3 + 3'h1; // @[Counter.scala 76:24]
  wire  releaseLast = _T_168 & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  respToL1Fire = hitReadBurst & _T_148; // @[Cache.scala 354:51]
  wire  _T_179 = _T_160 | _T_164; // @[Cache.scala 355:48]
  wire  _T_180 = (_T_160 | _T_164) & hitReadBurst; // @[Cache.scala 355:96]
  reg [2:0] value_4; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = value_4 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_3 = value_4 + 3'h1; // @[Counter.scala 76:24]
  wire  respToL1Last = _T_180 & wrap_wrap_1; // @[Counter.scala 118:{17,24}]
  wire [3:0] _T_184 = hit ? 4'h8 : 4'h0; // @[Cache.scala 364:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[Cache.scala 369:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[Cache.scala 369:33]
  wire [3:0] _T_191 = meta_dirty ? 4'h3 : 4'h1; // @[Cache.scala 371:42]
  wire [3:0] _T_192 = mmio ? 4'h5 : _T_191; // @[Cache.scala 371:21]
  wire [3:0] _GEN_20 = miss | mmio ? _T_192 : state; // @[Cache.scala 370:49 371:15 298:22]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : value_1; // @[Cache.scala 379:48 Counter.scala 76:15 60:40]
  wire  _T_203 = respToL1Fire & respToL1Last; // @[Cache.scala 380:71]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[Cache.scala 298:22 380:{88,96}]
  wire [3:0] _GEN_29 = _T_134 ? 4'h2 : state; // @[Cache.scala 383:50 384:13 298:22]
  wire [2:0] _GEN_30 = _T_134 ? addr_wordIndex : value_1; // @[Cache.scala 383:50 385:25 Counter.scala 60:40]
  wire [2:0] _GEN_31 = _T_86 ? 3'h0 : _GEN_0; // @[Cache.scala 392:{52,75}]
  wire  _T_210 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_210 ? 4'h7 : state; // @[Cache.scala 298:22 393:{46,54}]
  wire  _GEN_33 = _T_154 | afterFirstRead; // @[Cache.scala 389:33 390:24 340:31]
  wire [2:0] _GEN_34 = _T_154 ? _value_T_7 : value_1; // @[Cache.scala 389:33 Counter.scala 76:15 60:40]
  wire [2:0] _GEN_35 = _T_154 ? _GEN_31 : _GEN_0; // @[Cache.scala 389:33]
  wire [3:0] _GEN_36 = _T_154 ? _GEN_32 : state; // @[Cache.scala 298:22 389:33]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_134 ? _value_T_11 : value_2; // @[Cache.scala 398:32 Counter.scala 76:15 60:40]
  wire  _T_213 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_213 & _T_134 ? 4'h4 : state; // @[Cache.scala 298:22 399:{65,73}]
  wire [3:0] _GEN_39 = _T_154 ? 4'h1 : state; // @[Cache.scala 298:22 402:{53,61}]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[Cache.scala 298:22 403:{76,84}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[Cache.scala 357:18 298:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[Cache.scala 357:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : value_2; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[Cache.scala 357:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : value_1; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [2:0] _GEN_47 = 4'h2 == state ? _GEN_35 : _GEN_0; // @[Cache.scala 357:18]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[Cache.scala 357:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? value_2 : _GEN_43; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[Cache.scala 357:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[Cache.scala 357:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_53 = 4'h1 == state ? _GEN_0 : _GEN_47; // @[Cache.scala 357:18]
  wire [2:0] _GEN_54 = 4'h1 == state ? value_2 : _GEN_49; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[Cache.scala 357:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? _GEN_28 : _GEN_50; // @[Cache.scala 357:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[Cache.scala 357:18 340:31]
  wire [2:0] _GEN_58 = 4'h8 == state ? _GEN_0 : _GEN_53; // @[Cache.scala 357:18]
  wire [2:0] _GEN_59 = 4'h8 == state ? value_2 : _GEN_54; // @[Cache.scala 357:18 Counter.scala 60:40]
  wire [63:0] _T_222 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 406:67]
  wire [63:0] _T_223 = io_in_bits_req_wdata & _T_222; // @[BitUtils.scala 32:13]
  wire [63:0] _T_224 = ~_T_222; // @[BitUtils.scala 32:38]
  wire [63:0] _T_225 = io_mem_resp_bits_rdata & _T_224; // @[BitUtils.scala 32:36]
  wire [63:0] dataRefill = _T_223 | _T_225; // @[BitUtils.scala 32:25]
  wire  dataRefillWriteBus_req_valid = _T_156 & _T_154; // @[Cache.scala 408:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_210; // @[Cache.scala 416:61]
  wire  _T_246 = dataRefillWriteBus_req_valid & _T_7; // @[Cache.scala 426:59]
  wire [2:0] _T_248 = _T_210 ? 3'h6 : 3'h2; // @[Cache.scala 429:29]
  wire [63:0] _T_252 = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 432:31]
  wire [2:0] _T_255 = respToL1Last ? 3'h6 : 3'h2; // @[Cache.scala 437:29]
  wire [63:0] _GEN_76 = hitReadBurst & _T_111 ? _T_129 : _T_252; // @[Cache.scala 434:54 436:25 439:25]
  wire [3:0] _GEN_77 = hitReadBurst & _T_111 ? {{1'd0}, _T_255} : io_in_bits_req_cmd; // @[Cache.scala 434:54 437:23 440:23]
  wire [63:0] _GEN_78 = _T_87 | _T_86 ? _T_252 : _GEN_76; // @[Cache.scala 430:75 432:25]
  wire  _T_261 = state == 4'h7; // @[Cache.scala 450:48]
  wire  _T_274 = io_in_bits_req_cmd[0] & (hit | ~hit & state == 4'h7) | _T_246 | _T_203 & _T_111; // @[Cache.scala 450:161]
  wire  _T_280 = io_in_bits_req_cmd[0] | mmio ? _T_261 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 451:45]
  wire  _T_282 = probe ? 1'h0 : hit | _T_280; // @[Cache.scala 451:8]
  wire  _T_283 = io_in_bits_req_cmd[1] ? _T_274 : _T_282; // @[Cache.scala 449:37]
  wire  _T_289 = miss ? _T_160 : _T_111 & releaseLast; // @[Cache.scala 458:53]
  wire  _T_298 = hit | io_in_bits_req_cmd[0] ? io_out_valid : _T_261 & _GEN_12; // @[Cache.scala 459:8]
  Arbiter_10 metaWriteArb ( // @[Cache.scala 257:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_11 dataWriteArb ( // @[Cache.scala 258:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_160 & ~hitReadBurst & ~miss & ~probe; // @[Cache.scala 462:79]
  assign io_out_valid = io_in_valid & _T_283; // @[Cache.scala 449:31]
  assign io_out_bits_cmd = dataRefillWriteBus_req_valid & _T_7 ? {{1'd0}, _T_248} : _GEN_77; // @[Cache.scala 426:81 429:23]
  assign io_out_bits_rdata = dataRefillWriteBus_req_valid & _T_7 ? dataRefill : _GEN_78; // @[Cache.scala 426:81 428:25]
  assign io_isFinish = probe ? io_cohResp_valid & _T_289 : _T_298; // @[Cache.scala 458:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 310:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_116}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 413:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 413:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 423:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 423:23]
  assign io_mem_req_valid = _T_140 | _T_110 & state2 == 2'h2; // @[Cache.scala 333:48]
  assign io_mem_req_bits_addr = _T_140 ? raddr : waddr; // @[Cache.scala 328:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_128 | _T_126; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 332:21]
  assign io_cohResp_valid = state == 4'h0 & probe | _T_164; // @[Cache.scala 347:53]
  assign io_dataReadRespToL1 = hitReadBurst & _T_179; // @[Cache.scala 463:39]
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[Cache.scala 293:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 292:29 SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_210; // @[Cache.scala 416:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 261:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 415:32 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 287:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_98}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = _T_91 | _T_93; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 288:29 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _T_156 & _T_154; // @[Cache.scala 408:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = _T_223 | _T_225; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 407:32 SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      value <= _GEN_0;
    end else if (4'h5 == state) begin // @[Cache.scala 357:18]
      value <= _GEN_0;
    end else if (4'h6 == state) begin // @[Cache.scala 357:18]
      value <= _GEN_0;
    end else begin
      value <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 298:22]
      state <= 4'h0; // @[Cache.scala 298:22]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      if (probe) begin // @[Cache.scala 362:20]
        if (io_cohResp_valid) begin // @[Cache.scala 363:34]
          state <= _T_184; // @[Cache.scala 364:17]
        end
      end else if (hitReadBurst) begin // @[Cache.scala 367:50]
        state <= 4'h8; // @[Cache.scala 368:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
        state <= _GEN_56;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      if (probe) begin // @[Cache.scala 362:20]
        if (io_cohResp_valid) begin // @[Cache.scala 363:34]
          value_1 <= addr_wordIndex; // @[Cache.scala 365:29]
        end
      end else if (hitReadBurst) begin // @[Cache.scala 367:50]
        value_1 <= _value_T_5; // @[Cache.scala 369:27]
      end
    end else if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
        value_1 <= _GEN_55;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 308:23]
      state2 <= 2'h0; // @[Cache.scala 308:23]
    end else if (2'h0 == state2) begin // @[Cache.scala 315:19]
      if (_T_131) begin // @[Cache.scala 316:53]
        state2 <= 2'h1; // @[Cache.scala 316:62]
      end
    end else if (2'h1 == state2) begin // @[Cache.scala 315:19]
      state2 <= 2'h2; // @[Cache.scala 317:35]
    end else if (2'h2 == state2) begin // @[Cache.scala 315:19]
      state2 <= _GEN_8;
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 16:23]
    end
    if (_T_118) begin // @[Reg.scala 16:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Cache.scala 340:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 340:31]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      afterFirstRead <= 1'h0; // @[Cache.scala 359:22]
    end else if (!(4'h5 == state)) begin // @[Cache.scala 357:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 357:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (4'h0 == state) begin // @[Cache.scala 357:18]
      alreadyOutFire <= 1'h0; // @[Cache.scala 360:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_159) begin // @[Reg.scala 16:19]
      if (mmio) begin // @[Cache.scala 343:39]
        inRdataRegDemand <= 64'h0;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_3 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_168) begin // @[Counter.scala 118:17]
      value_3 <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_4 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_180) begin // @[Counter.scala 118:17]
      value_4 <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:268 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 268:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 268:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:465 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 465:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 465:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:466 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 466:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 466:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  value_3 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  value_4 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_5(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [8:0]  io_rreq_bits_setIdx,
  output [16:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [16:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [16:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [16:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [16:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  reg  REG; // @[SRAMTemplate.scala 80:30]
  reg [8:0] value; // @[Counter.scala 60:40]
  wire  wrap_wrap = value == 9'h1ff; // @[Counter.scala 72:24]
  wire [8:0] _wrap_value_T_1 = value + 9'h1; // @[Counter.scala 76:24]
  wire  wrap = REG & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = wrap ? 1'h0 : REG; // @[SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  wire  _T = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = REG ? value : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [18:0] _T_1 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = REG ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [18:0] _WIRE_2 = array_RW0_rdata_0;
  wire [18:0] _WIRE_3 = array_RW0_rdata_1;
  wire [18:0] _WIRE_4 = array_RW0_rdata_2;
  wire [18:0] _WIRE_5 = array_RW0_rdata_3;
  array_2 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~REG & _T; // @[SRAMTemplate.scala 101:33]
  assign io_rresp_data_0_tag = _WIRE_2[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_valid = _WIRE_2[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_dirty = _WIRE_2[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_tag = _WIRE_3[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_valid = _WIRE_3[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_dirty = _WIRE_3[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_tag = _WIRE_4[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_valid = _WIRE_4[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_dirty = _WIRE_4[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_tag = _WIRE_5[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_valid = _WIRE_5[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_dirty = _WIRE_5[0]; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | wen;
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[Counter.scala 60:40]
      value <= 9'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      value <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_12(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [8:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [8:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter_4(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [8:0]  io_r0_req_bits_setIdx,
  output [16:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [16:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [16:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [16:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [16:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [16:0] r_0_tag; // @[Reg.scala 27:20]
  reg  r_0_valid; // @[Reg.scala 27:20]
  reg  r_0_dirty; // @[Reg.scala 27:20]
  reg [16:0] r_1_tag; // @[Reg.scala 27:20]
  reg  r_1_valid; // @[Reg.scala 27:20]
  reg  r_1_dirty; // @[Reg.scala 27:20]
  reg [16:0] r_2_tag; // @[Reg.scala 27:20]
  reg  r_2_valid; // @[Reg.scala 27:20]
  reg  r_2_dirty; // @[Reg.scala 27:20]
  reg [16:0] r_3_tag; // @[Reg.scala 27:20]
  reg  r_3_valid; // @[Reg.scala 27:20]
  reg  r_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_5 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_12 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_tag = REG ? ram_io_rresp_data_0_tag : r_0_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_valid = REG ? ram_io_rresp_data_0_valid : r_0_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_dirty = REG ? ram_io_rresp_data_0_dirty : r_0_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_tag = REG ? ram_io_rresp_data_1_tag : r_1_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_valid = REG ? ram_io_rresp_data_1_valid : r_1_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_dirty = REG ? ram_io_rresp_data_1_dirty : r_1_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_tag = REG ? ram_io_rresp_data_2_tag : r_2_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_valid = REG ? ram_io_rresp_data_2_valid : r_2_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_dirty = REG ? ram_io_rresp_data_2_dirty : r_2_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_tag = REG ? ram_io_rresp_data_3_tag : r_3_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_valid = REG ? ram_io_rresp_data_3_valid : r_3_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_dirty = REG ? ram_io_rresp_data_3_dirty : r_3_dirty; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_0_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_tag <= ram_io_rresp_data_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_valid <= ram_io_rresp_data_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_dirty <= ram_io_rresp_data_0_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_tag <= ram_io_rresp_data_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_valid <= ram_io_rresp_data_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_dirty <= ram_io_rresp_data_1_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_tag <= ram_io_rresp_data_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_valid <= ram_io_rresp_data_2_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_dirty <= ram_io_rresp_data_2_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_tag <= ram_io_rresp_data_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_valid <= ram_io_rresp_data_3_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_dirty <= ram_io_rresp_data_3_dirty; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_0_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  r_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_tag = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_2_tag = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  r_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_3_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  r_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_6(
  input         clock,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [11:0] io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [11:0] io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire [11:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  wire  realRen = io_rreq_valid & ~io_wreq_valid; // @[SRAMTemplate.scala 89:38]
  array_3 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 101:53]
  assign io_rresp_data_0_data = array_RW0_rdata_0; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_data = array_RW0_rdata_1; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_data = array_RW0_rdata_2; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_data = array_RW0_rdata_3; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = io_wreq_bits_waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = io_wreq_bits_waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = io_wreq_bits_waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = io_wreq_bits_waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | io_wreq_valid;
  assign array_RW0_wmode = io_wreq_valid; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx;
endmodule
module Arbiter_13(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module SRAMTemplateWithArbiter_5(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [11:0] io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [11:0] io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [11:0] io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r__0_data; // @[Reg.scala 27:20]
  reg [63:0] r__1_data; // @[Reg.scala 27:20]
  reg [63:0] r__2_data; // @[Reg.scala 27:20]
  reg [63:0] r__3_data; // @[Reg.scala 27:20]
  reg  REG_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r_1_0_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_1_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_2_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_6 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_13 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_data = REG ? ram_io_rresp_data_0_data : r__0_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_data = REG ? ram_io_rresp_data_1_data : r__1_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_data = REG ? ram_io_rresp_data_2_data : r__2_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_data = REG ? ram_io_rresp_data_3_data : r__3_data; // @[Hold.scala 23:48]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r1_resp_data_0_data = REG_1 ? ram_io_rresp_data_0_data : r_1_0_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_1_data = REG_1 ? ram_io_rresp_data_1_data : r_1_1_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_2_data = REG_1 ? ram_io_rresp_data_2_data : r_1_2_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_3_data = REG_1 ? ram_io_rresp_data_3_data : r_1_3_data; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r__0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
    REG_1 <= io_r1_req_ready & io_r1_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_1_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r__0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r__1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  r__2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  r__3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  r_1_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  r_1_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 484:18]
  wire  s1_io_in_valid; // @[Cache.scala 484:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 484:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 484:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 484:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 484:18]
  wire  s1_io_out_ready; // @[Cache.scala 484:18]
  wire  s1_io_out_valid; // @[Cache.scala 484:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 484:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 484:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 484:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 484:18]
  wire [8:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [16:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 484:18]
  wire [16:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 484:18]
  wire [16:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 484:18]
  wire [16:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 484:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 484:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 484:18]
  wire [11:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 484:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 484:18]
  wire  s2_clock; // @[Cache.scala 485:18]
  wire  s2_reset; // @[Cache.scala 485:18]
  wire  s2_io_in_ready; // @[Cache.scala 485:18]
  wire  s2_io_in_valid; // @[Cache.scala 485:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 485:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 485:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 485:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 485:18]
  wire  s2_io_out_ready; // @[Cache.scala 485:18]
  wire  s2_io_out_valid; // @[Cache.scala 485:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 485:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 485:18]
  wire [16:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 485:18]
  wire [16:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 485:18]
  wire [16:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 485:18]
  wire [16:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 485:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 485:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 485:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 485:18]
  wire [16:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 485:18]
  wire [16:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 485:18]
  wire [16:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 485:18]
  wire [16:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 485:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 485:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 485:18]
  wire [8:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 485:18]
  wire [16:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 485:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 485:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 485:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 485:18]
  wire [11:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 485:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 485:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 485:18]
  wire  s3_clock; // @[Cache.scala 486:18]
  wire  s3_reset; // @[Cache.scala 486:18]
  wire  s3_io_in_ready; // @[Cache.scala 486:18]
  wire  s3_io_in_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 486:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 486:18]
  wire [16:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 486:18]
  wire [16:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 486:18]
  wire [16:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 486:18]
  wire [16:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 486:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 486:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 486:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 486:18]
  wire  s3_io_out_valid; // @[Cache.scala 486:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_isFinish; // @[Cache.scala 486:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 486:18]
  wire [11:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 486:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 486:18]
  wire [11:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 486:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 486:18]
  wire [8:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 486:18]
  wire [16:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 486:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 486:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 486:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 486:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 486:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 486:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 486:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 486:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 486:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 486:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 486:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 486:18]
  wire  metaArray_clock; // @[Cache.scala 487:25]
  wire  metaArray_reset; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 487:25]
  wire [8:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 487:25]
  wire [16:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 487:25]
  wire [16:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 487:25]
  wire [16:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 487:25]
  wire [16:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 487:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 487:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 487:25]
  wire [8:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 487:25]
  wire [16:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 487:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 487:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 487:25]
  wire  dataArray_clock; // @[Cache.scala 488:25]
  wire  dataArray_reset; // @[Cache.scala 488:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 488:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 488:25]
  wire [11:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 488:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 488:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 488:25]
  wire [11:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 488:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 488:25]
  wire [11:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 488:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 488:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 488:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 497:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 497:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 497:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 497:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 497:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 497:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 497:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 497:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 497:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 497:19]
  wire  arb_io_out_ready; // @[Cache.scala 497:19]
  wire  arb_io_out_valid; // @[Cache.scala 497:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 497:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 497:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 497:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 497:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 497:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_req_addr; // @[Reg.scala 15:16]
  reg [3:0] r_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_req_wdata; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_5 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [3:0] r_1_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_1_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_1_req_wdata; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_0_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_0_dirty; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_1_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_1_dirty; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_2_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_2_dirty; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_3_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_3_data; // @[Reg.scala 15:16]
  reg  r_1_hit; // @[Reg.scala 15:16]
  reg [3:0] r_1_waymask; // @[Reg.scala 15:16]
  reg  r_1_mmio; // @[Reg.scala 15:16]
  reg  r_1_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] r_1_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] r_1_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_11 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  CacheStage1_2 s1 ( // @[Cache.scala 484:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2_2 s2 ( // @[Cache.scala 485:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3_2 s3 ( // @[Cache.scala 486:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  SRAMTemplateWithArbiter_4 metaArray ( // @[Cache.scala 487:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_5 dataArray ( // @[Cache.scala 488:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 497:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 498:28]
  assign io_in_resp_valid = s3_io_out_valid & _T_11 ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 514:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 508:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 508:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 510:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 510:14]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 500:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 500:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 500:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 500:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 500:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 532:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 532:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 533:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 533:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = r_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = r_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = r_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = r_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 539:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 539:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 540:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 542:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 542:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 541:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 541:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = r_1_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = r_1_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = r_1_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = r_1_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = r_1_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = r_1_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = r_1_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = r_1_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = r_1_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = r_1_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = r_1_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = r_1_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = r_1_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = r_1_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = r_1_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = r_1_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = r_1_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = r_1_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = r_1_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = r_1_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = r_1_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = r_1_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 534:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 534:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 510:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 510:14]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 532:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 532:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 536:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 536:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 533:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 533:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 534:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 534:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 537:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 537:18]
  assign arb_io_in_0_valid = 1'h0; // @[Cache.scala 522:24]
  assign arb_io_in_0_bits_addr = 32'h0; // @[Cache.scala 519:19 SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_size = 3'h0; // @[Cache.scala 519:19 SimpleBus.scala 66:15]
  assign arb_io_in_0_bits_cmd = 4'h0; // @[Cache.scala 519:19 SimpleBus.scala 65:14]
  assign arb_io_in_0_bits_wmask = 8'h0; // @[Cache.scala 519:19 SimpleBus.scala 68:16]
  assign arb_io_in_0_bits_wdata = 64'h0; // @[Cache.scala 519:19 SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 498:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 498:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 500:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_cmd <= s1_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wmask <= s1_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wdata <= s1_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_1 <= _GEN_9;
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_cmd <= s2_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wmask <= s2_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wdata <= s2_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_hit <= s2_io_out_bits_hit; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_req_cmd = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  r_req_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  r_req_wdata = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_req_addr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_req_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_req_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_req_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_metas_0_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  r_1_metas_0_dirty = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_1_metas_1_tag = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  r_1_metas_1_dirty = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_1_metas_2_tag = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  r_1_metas_2_dirty = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_metas_3_tag = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_metas_3_dirty = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  r_1_datas_0_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  r_1_datas_1_data = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  r_1_datas_2_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  r_1_datas_3_data = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  r_1_hit = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_1_waymask = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  r_1_mmio = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_1_isForwardData = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  r_1_forwardData_data_data = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  r_1_forwardData_waymask = _RAND_27[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusAddressMapper(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [3:0]  io_out_req_bits_cmd,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
  assign io_in_req_ready = io_out_req_ready; // @[AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = {4'h8,io_in_req_bits_addr[27:0]}; // @[Cat.scala 30:58]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [2:0]  io_out_awprot,
  output        io_out_awid,
  output        io_out_awuser,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  output        io_out_awlock,
  output [3:0]  io_out_awcache,
  output [3:0]  io_out_awqos,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output        io_out_wlast,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [2:0]  io_out_arprot,
  output        io_out_arid,
  output        io_out_aruser,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_arlock,
  output [3:0]  io_out_arcache,
  output [3:0]  io_out_arqos,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_13 & _T_17 & io_out_wlast | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_28 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_36 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awprot = io_out_arprot; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awuser = io_out_aruser; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_awlock = io_out_arlock; // @[ToAXI4.scala 182:6]
  assign io_out_awcache = io_out_arcache; // @[ToAXI4.scala 182:6]
  assign io_out_awqos = io_out_arqos; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:54]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arprot = 3'h1; // @[ToAXI4.scala 159:12]
  assign io_out_arid = 1'h0; // @[ToAXI4.scala 168:24]
  assign io_out_aruser = 1'h0; // @[ToAXI4.scala 176:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_arsize = 3'h3; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h2; // @[ToAXI4.scala 171:24]
  assign io_out_arlock = 1'h0; // @[ToAXI4.scala 173:24]
  assign io_out_arcache = 4'h0; // @[ToAXI4.scala 174:24]
  assign io_out_arqos = 4'h0; // @[ToAXI4.scala 175:24]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin // @[Reg.scala 16:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [2:0]  io_out_2_req_bits_size,
  output [3:0]  io_out_2_req_bits_cmd,
  output [7:0]  io_out_2_req_bits_wmask,
  output [63:0] io_out_2_req_bits_wdata,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [3:0]  io_out_2_resp_bits_cmd,
  input  [63:0] io_out_2_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h38000000 & io_in_req_bits_addr < 32'h38010000; // @[Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h3c000000 & io_in_req_bits_addr < 32'h40000000; // @[Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40600000 & io_in_req_bits_addr < 32'h41600000; // @[Crossbar.scala 37:34]
  wire [2:0] _enc_T = outMatchVec_2 ? 3'h4 : 3'h0; // @[Mux.scala 47:69]
  wire [2:0] _enc_T_1 = outMatchVec_1 ? 3'h2 : _enc_T; // @[Mux.scala 47:69]
  wire [2:0] enc = outMatchVec_0 ? 3'h1 : _enc_T_1; // @[Mux.scala 47:69]
  wire  outSelVec_0 = enc[0]; // @[OneHot.scala 83:30]
  wire  outSelVec_1 = enc[1]; // @[OneHot.scala 83:30]
  wire  outSelVec_2 = enc[2]; // @[OneHot.scala 83:30]
  wire  _T_12 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_13 = state == 2'h0; // @[Crossbar.scala 41:66]
  wire  _T_14 = _T_12 & state == 2'h0; // @[Crossbar.scala 41:57]
  reg  outSelRespVec_0; // @[Reg.scala 27:20]
  reg  outSelRespVec_1; // @[Reg.scala 27:20]
  reg  outSelRespVec_2; // @[Reg.scala 27:20]
  wire [2:0] _T_15 = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_T_15); // @[Crossbar.scala 42:40]
  wire [1:0] _GEN_5 = io_in_resp_valid ? 2'h0 : state; // @[Crossbar.scala 32:22 56:{44,52}]
  wire  _T_37 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 & io_out_2_req_ready; // @[Mux.scala 27:72]
  wire  _T_61 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid | outSelRespVec_2 &
    io_out_2_resp_valid; // @[Mux.scala 27:72]
  wire [63:0] _T_64 = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_65 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_66 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_67 = _T_64 | _T_65; // @[Mux.scala 27:72]
  wire [3:0] _T_69 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_70 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_71 = outSelRespVec_2 ? io_out_2_resp_bits_cmd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_72 = _T_69 | _T_70; // @[Mux.scala 27:72]
  assign io_in_req_ready = _T_37 | reqInvalidAddr; // @[Crossbar.scala 61:64]
  assign io_in_resp_valid = _T_61 | state == 2'h2; // @[Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _T_72 | _T_71; // @[Mux.scala 27:72]
  assign io_in_resp_bits_rdata = _T_67 | _T_66; // @[Mux.scala 27:72]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _T_13; // @[Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & state == 2'h1; // @[Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _T_13; // @[Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & state == 2'h1; // @[Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _T_13; // @[Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 64:24]
  assign io_out_2_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & state == 2'h1; // @[Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 32:22]
      state <= 2'h0; // @[Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[Crossbar.scala 54:29]
        state <= 2'h2; // @[Crossbar.scala 54:37]
      end else if (_T_12) begin // @[Crossbar.scala 53:31]
        state <= 2'h1; // @[Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[Crossbar.scala 51:18]
      state <= _GEN_5;
    end else if (2'h2 == state) begin // @[Crossbar.scala 51:18]
      state <= _GEN_5;
    end
    if (reset) begin // @[Reg.scala 27:20]
      outSelRespVec_0 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_14) begin // @[Reg.scala 28:19]
      outSelRespVec_0 <= outSelVec_0; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      outSelRespVec_1 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_14) begin // @[Reg.scala 28:19]
      outSelRespVec_1 <= outSelVec_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      outSelRespVec_2 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_14) begin // @[Reg.scala 28:19]
      outSelRespVec_2 <= outSelVec_2; // @[Reg.scala 28:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~reqInvalidAddr | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~reqInvalidAddr | reset)) begin
          $fatal; // @[Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [2:0]  io_out_awprot,
  output        io_out_awid,
  output        io_out_awuser,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  output        io_out_awlock,
  output [3:0]  io_out_awcache,
  output [3:0]  io_out_awqos,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_wlast,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [2:0]  io_out_arprot,
  output        io_out_arid,
  output        io_out_aruser,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_arlock,
  output [3:0]  io_out_arcache,
  output [3:0]  io_out_arqos,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_13 & _T_17 & io_out_wlast | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_28 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_36 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awprot = io_out_arprot; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awuser = io_out_aruser; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_awlock = io_out_arlock; // @[ToAXI4.scala 182:6]
  assign io_out_awcache = io_out_arcache; // @[ToAXI4.scala 182:6]
  assign io_out_awqos = io_out_arqos; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:54]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arprot = 3'h1; // @[ToAXI4.scala 159:12]
  assign io_out_arid = 1'h0; // @[ToAXI4.scala 168:24]
  assign io_out_aruser = 1'h0; // @[ToAXI4.scala 176:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_arsize = io_in_req_bits_size; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h1; // @[ToAXI4.scala 171:24]
  assign io_out_arlock = 1'h0; // @[ToAXI4.scala 173:24]
  assign io_out_arcache = 4'h0; // @[ToAXI4.scala 174:24]
  assign io_out_arqos = 4'h0; // @[ToAXI4.scala 175:24]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin // @[Reg.scala 16:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  output        io__extra_mtip,
  output        io__extra_msip,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _T_9 = io__in_wstrb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_11 = io__in_wstrb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_13 = io__in_wstrb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_15 = io__in_wstrb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_17 = io__in_wstrb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_19 = io__in_wstrb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_21 = io__in_wstrb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_23 = io__in_wstrb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] fullMask = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 30:58]
  wire  _T_24 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_25 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_25 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_25 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  reg [63:0] mtime; // @[AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[AXI4CLINT.scala 34:21]
  reg [15:0] freq; // @[AXI4CLINT.scala 37:21]
  reg [15:0] inc; // @[AXI4CLINT.scala 38:20]
  reg [15:0] cnt; // @[AXI4CLINT.scala 40:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[AXI4CLINT.scala 41:21]
  wire  tick = nextCnt == freq; // @[AXI4CLINT.scala 43:23]
  wire [63:0] _GEN_14 = {{48'd0}, inc}; // @[AXI4CLINT.scala 44:32]
  wire [63:0] _T_49 = mtime + _GEN_14; // @[AXI4CLINT.scala 44:32]
  wire  _T_78 = 16'h0 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_79 = 16'h8000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_80 = 16'hbff8 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_81 = 16'h8008 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_82 = 16'h4000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_83 = _T_78 ? msip : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_84 = _T_79 ? freq : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_85 = _T_80 ? mtime : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_86 = _T_81 ? inc : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_87 = _T_82 ? mtimecmp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_15 = {{48'd0}, _T_84}; // @[Mux.scala 27:72]
  wire [63:0] _T_88 = _T_83 | _GEN_15; // @[Mux.scala 27:72]
  wire [63:0] _T_89 = _T_88 | _T_85; // @[Mux.scala 27:72]
  wire [63:0] _GEN_16 = {{48'd0}, _T_86}; // @[Mux.scala 27:72]
  wire [63:0] _T_90 = _T_89 | _GEN_16; // @[Mux.scala 27:72]
  wire [63:0] _T_94 = io__in_wdata & fullMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_95 = ~fullMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_96 = msip & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_97 = _T_94 | _T_96; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_17 = {{48'd0}, freq}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_102 = _GEN_17 & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_103 = _T_94 | _T_102; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_10 = _T_42 & io__in_awaddr[15:0] == 16'h8000 ? _T_103 : {{48'd0}, freq}; // @[RegMap.scala 32:{48,52} AXI4CLINT.scala 37:21]
  wire [63:0] _T_108 = mtime & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_109 = _T_94 | _T_108; // @[BitUtils.scala 32:25]
  wire [63:0] _T_114 = _GEN_14 & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_115 = _T_94 | _T_114; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_12 = _T_42 & io__in_awaddr[15:0] == 16'h8008 ? _T_115 : {{48'd0}, inc}; // @[RegMap.scala 32:{48,52} AXI4CLINT.scala 38:20]
  wire [63:0] _T_120 = mtimecmp & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_121 = _T_94 | _T_120; // @[BitUtils.scala 32:25]
  reg  REG_3; // @[AXI4CLINT.scala 64:31]
  reg  REG_4; // @[AXI4CLINT.scala 65:31]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io__in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io__in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = _T_90 | _T_87; // @[Mux.scala 27:72]
  assign io__extra_mtip = REG_3; // @[AXI4CLINT.scala 64:21]
  assign io__extra_msip = REG_4; // @[AXI4CLINT.scala 65:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    if (reset) begin // @[AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[AXI4CLINT.scala 32:22]
    end else if (_T_42 & io__in_awaddr[15:0] == 16'hbff8) begin // @[RegMap.scala 32:48]
      mtime <= _T_109; // @[RegMap.scala 32:52]
    end else if (tick) begin // @[AXI4CLINT.scala 44:15]
      mtime <= _T_49; // @[AXI4CLINT.scala 44:23]
    end
    if (reset) begin // @[AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[AXI4CLINT.scala 33:25]
    end else if (_T_42 & io__in_awaddr[15:0] == 16'h4000) begin // @[RegMap.scala 32:48]
      mtimecmp <= _T_121; // @[RegMap.scala 32:52]
    end
    if (reset) begin // @[AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[AXI4CLINT.scala 34:21]
    end else if (_T_42 & io__in_awaddr[15:0] == 16'h0) begin // @[RegMap.scala 32:48]
      msip <= _T_97; // @[RegMap.scala 32:52]
    end
    if (reset) begin // @[AXI4CLINT.scala 37:21]
      freq <= 16'h64; // @[AXI4CLINT.scala 37:21]
    end else begin
      freq <= _GEN_10[15:0];
    end
    if (reset) begin // @[AXI4CLINT.scala 38:20]
      inc <= 16'h1; // @[AXI4CLINT.scala 38:20]
    end else begin
      inc <= _GEN_12[15:0];
    end
    if (reset) begin // @[AXI4CLINT.scala 40:20]
      cnt <= 16'h0; // @[AXI4CLINT.scala 40:20]
    end else if (nextCnt < freq) begin // @[AXI4CLINT.scala 42:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    REG_3 <= mtime >= mtimecmp; // @[AXI4CLINT.scala 64:38]
    REG_4 <= msip != 64'h0; // @[AXI4CLINT.scala 65:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  freq = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inc = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  REG_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_4 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBus2AXI4Converter_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[ToAXI4.scala 151:20]
  wire  _T_8 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_8 | awAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_12 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_8 & _T_12 | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _GEN_2 = _T_12 | wAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_18 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_23 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_26 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_31 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_31 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_26 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_26 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_23; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_18) begin // @[Reg.scala 16:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(toAXI4Lite | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(toAXI4Lite | reset)) begin
          $fatal; // @[ToAXI4.scala 153:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  input  [2:0]  io__extra_intrVec,
  output        io__extra_meip_0,
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _T_24 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_25 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_25 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_25 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  reg [31:0] priority_0; // @[AXI4PLIC.scala 37:39]
  reg [31:0] priority_1; // @[AXI4PLIC.scala 37:39]
  reg [31:0] priority_2; // @[AXI4PLIC.scala 37:39]
  reg  pending_0_1; // @[AXI4PLIC.scala 43:46]
  reg  pending_0_2; // @[AXI4PLIC.scala 43:46]
  reg  pending_0_3; // @[AXI4PLIC.scala 43:46]
  wire [31:0] _T_45 = {16'h0,8'h0,4'h0,pending_0_3,pending_0_2,pending_0_1,1'h0}; // @[Cat.scala 30:58]
  reg [31:0] enable_0_0; // @[AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[AXI4PLIC.scala 53:40]
  reg  inHandle_1; // @[AXI4PLIC.scala 58:25]
  reg  inHandle_2; // @[AXI4PLIC.scala 58:25]
  reg  inHandle_3; // @[AXI4PLIC.scala 58:25]
  reg [31:0] claimCompletion_0; // @[AXI4PLIC.scala 64:46]
  wire  _GEN_13 = _T_25 & io__in_araddr[25:0] == 26'h200004 ? 2'h1 == claimCompletion_0[1:0] | inHandle_1 :
    inHandle_1; // @[AXI4PLIC.scala 58:25 68:59]
  wire  _GEN_14 = _T_25 & io__in_araddr[25:0] == 26'h200004 ? 2'h2 == claimCompletion_0[1:0] | inHandle_2 :
    inHandle_2; // @[AXI4PLIC.scala 58:25 68:59]
  wire  _GEN_15 = _T_25 & io__in_araddr[25:0] == 26'h200004 ? 2'h3 == claimCompletion_0[1:0] | inHandle_3 :
    inHandle_3; // @[AXI4PLIC.scala 58:25 68:59]
  wire  _GEN_16 = io__extra_intrVec[0] | pending_0_1; // @[AXI4PLIC.scala 75:{17,45} 43:46]
  wire  _GEN_18 = io__extra_intrVec[1] | pending_0_2; // @[AXI4PLIC.scala 75:{17,45} 43:46]
  wire  _GEN_20 = io__extra_intrVec[2] | pending_0_3; // @[AXI4PLIC.scala 75:{17,45} 43:46]
  wire [31:0] _T_54 = _T_45 & enable_0_0; // @[AXI4PLIC.scala 81:31]
  wire [4:0] _T_88 = _T_54[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  wire [4:0] _T_89 = _T_54[29] ? 5'h1d : _T_88; // @[Mux.scala 47:69]
  wire [4:0] _T_90 = _T_54[28] ? 5'h1c : _T_89; // @[Mux.scala 47:69]
  wire [4:0] _T_91 = _T_54[27] ? 5'h1b : _T_90; // @[Mux.scala 47:69]
  wire [4:0] _T_92 = _T_54[26] ? 5'h1a : _T_91; // @[Mux.scala 47:69]
  wire [4:0] _T_93 = _T_54[25] ? 5'h19 : _T_92; // @[Mux.scala 47:69]
  wire [4:0] _T_94 = _T_54[24] ? 5'h18 : _T_93; // @[Mux.scala 47:69]
  wire [4:0] _T_95 = _T_54[23] ? 5'h17 : _T_94; // @[Mux.scala 47:69]
  wire [4:0] _T_96 = _T_54[22] ? 5'h16 : _T_95; // @[Mux.scala 47:69]
  wire [4:0] _T_97 = _T_54[21] ? 5'h15 : _T_96; // @[Mux.scala 47:69]
  wire [4:0] _T_98 = _T_54[20] ? 5'h14 : _T_97; // @[Mux.scala 47:69]
  wire [4:0] _T_99 = _T_54[19] ? 5'h13 : _T_98; // @[Mux.scala 47:69]
  wire [4:0] _T_100 = _T_54[18] ? 5'h12 : _T_99; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = _T_54[17] ? 5'h11 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = _T_54[16] ? 5'h10 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = _T_54[15] ? 5'hf : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = _T_54[14] ? 5'he : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = _T_54[13] ? 5'hd : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = _T_54[12] ? 5'hc : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = _T_54[11] ? 5'hb : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = _T_54[10] ? 5'ha : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = _T_54[9] ? 5'h9 : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = _T_54[8] ? 5'h8 : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = _T_54[7] ? 5'h7 : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = _T_54[6] ? 5'h6 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = _T_54[5] ? 5'h5 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = _T_54[4] ? 5'h4 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = _T_54[3] ? 5'h3 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = _T_54[2] ? 5'h2 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = _T_54[1] ? 5'h1 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = _T_54[0] ? 5'h0 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = _T_54 == 32'h0 ? 5'h0 : _T_118; // @[AXI4PLIC.scala 82:13]
  wire [7:0] _T_124 = io__in_wstrb >> io__in_awaddr[2:0]; // @[AXI4PLIC.scala 89:78]
  wire [7:0] _T_134 = _T_124[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_136 = _T_124[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_138 = _T_124[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_140 = _T_124[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_142 = _T_124[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_144 = _T_124[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_146 = _T_124[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_148 = _T_124[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_149 = {_T_148,_T_146,_T_144,_T_142,_T_140,_T_138,_T_136,_T_134}; // @[Cat.scala 30:58]
  wire  _T_150 = 26'hc == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_151 = 26'h1000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_152 = 26'h2000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_153 = 26'h8 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_154 = 26'h200004 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_155 = 26'h4 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_156 = 26'h200000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_157 = _T_150 ? priority_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_158 = _T_151 ? _T_45 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_159 = _T_152 ? enable_0_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_160 = _T_153 ? priority_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_161 = _T_154 ? claimCompletion_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_162 = _T_155 ? priority_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_163 = _T_156 ? threshold_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_164 = _T_157 | _T_158; // @[Mux.scala 27:72]
  wire [31:0] _T_165 = _T_164 | _T_159; // @[Mux.scala 27:72]
  wire [31:0] _T_166 = _T_165 | _T_160; // @[Mux.scala 27:72]
  wire [31:0] _T_167 = _T_166 | _T_161; // @[Mux.scala 27:72]
  wire [31:0] _T_168 = _T_167 | _T_162; // @[Mux.scala 27:72]
  wire [31:0] rdata = _T_168 | _T_163; // @[Mux.scala 27:72]
  wire [63:0] _T_172 = io__in_wdata & _T_149; // @[BitUtils.scala 32:13]
  wire [63:0] _T_173 = ~_T_149; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_40 = {{32'd0}, priority_2}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_174 = _GEN_40 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_175 = _T_172 | _T_174; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_22 = _T_42 & io__in_awaddr[25:0] == 26'hc ? _T_175 : {{32'd0}, priority_2}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 37:39]
  wire [63:0] _GEN_41 = {{32'd0}, enable_0_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_180 = _GEN_41 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_181 = _T_172 | _T_180; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_23 = _T_42 & io__in_awaddr[25:0] == 26'h2000 ? _T_181 : {{32'd0}, enable_0_0}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 48:64]
  wire [63:0] _GEN_42 = {{32'd0}, priority_1}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_186 = _GEN_42 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_187 = _T_172 | _T_186; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_24 = _T_42 & io__in_awaddr[25:0] == 26'h8 ? _T_187 : {{32'd0}, priority_1}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 37:39]
  wire [63:0] _GEN_43 = {{32'd0}, claimCompletion_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_192 = _GEN_43 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_193 = _T_172 | _T_192; // @[BitUtils.scala 32:25]
  wire [4:0] _GEN_33 = _T_42 & io__in_awaddr[25:0] == 26'h200004 ? 5'h0 : _T_119; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 82:7]
  wire [63:0] _GEN_44 = {{32'd0}, priority_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_200 = _GEN_44 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_201 = _T_172 | _T_200; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_34 = _T_42 & io__in_awaddr[25:0] == 26'h4 ? _T_201 : {{32'd0}, priority_0}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 37:39]
  wire [63:0] _GEN_45 = {{32'd0}, threshold_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_206 = _GEN_45 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_207 = _T_172 | _T_206; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_35 = _T_42 & io__in_awaddr[25:0] == 26'h200000 ? _T_207 : {{32'd0}, threshold_0}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 53:40]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io__in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io__in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = {rdata,rdata}; // @[Cat.scala 30:58]
  assign io__extra_meip_0 = claimCompletion_0 != 32'h0; // @[AXI4PLIC.scala 93:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    priority_0 <= _GEN_34[31:0];
    priority_1 <= _GEN_24[31:0];
    priority_2 <= _GEN_22[31:0];
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_1 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_1) begin // @[AXI4PLIC.scala 76:25]
      pending_0_1 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_1 <= _GEN_16;
    end
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_2 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_2) begin // @[AXI4PLIC.scala 76:25]
      pending_0_2 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_2 <= _GEN_18;
    end
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_3 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_3) begin // @[AXI4PLIC.scala 76:25]
      pending_0_3 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_3 <= _GEN_20;
    end
    if (reset) begin // @[AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[AXI4PLIC.scala 48:64]
    end else begin
      enable_0_0 <= _GEN_23[31:0];
    end
    threshold_0 <= _GEN_35[31:0];
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_1 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_42 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (2'h1 == _T_193[1:0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_1 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_1 <= _GEN_13;
      end
    end else begin
      inHandle_1 <= _GEN_13;
    end
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_2 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_42 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (2'h2 == _T_193[1:0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_2 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_2 <= _GEN_14;
      end
    end else begin
      inHandle_2 <= _GEN_14;
    end
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_3 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_42 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (2'h3 == _T_193[1:0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_3 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_3 <= _GEN_15;
      end
    end else begin
      inHandle_3 <= _GEN_15;
    end
    claimCompletion_0 <= {{27'd0}, _GEN_33};
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  priority_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  priority_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  pending_0_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pending_0_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pending_0_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  enable_0_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  threshold_0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  inHandle_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inHandle_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inHandle_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  claimCompletion_0 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_awready,
  output        io_mem_awvalid,
  output [31:0] io_mem_awaddr,
  output [2:0]  io_mem_awprot,
  output        io_mem_awid,
  output        io_mem_awuser,
  output [7:0]  io_mem_awlen,
  output [2:0]  io_mem_awsize,
  output [1:0]  io_mem_awburst,
  output        io_mem_awlock,
  output [3:0]  io_mem_awcache,
  output [3:0]  io_mem_awqos,
  input         io_mem_wready,
  output        io_mem_wvalid,
  output [63:0] io_mem_wdata,
  output [7:0]  io_mem_wstrb,
  output        io_mem_wlast,
  output        io_mem_bready,
  input         io_mem_bvalid,
  input  [1:0]  io_mem_bresp,
  input         io_mem_bid,
  input         io_mem_buser,
  input         io_mem_arready,
  output        io_mem_arvalid,
  output [31:0] io_mem_araddr,
  output [2:0]  io_mem_arprot,
  output        io_mem_arid,
  output        io_mem_aruser,
  output [7:0]  io_mem_arlen,
  output [2:0]  io_mem_arsize,
  output [1:0]  io_mem_arburst,
  output        io_mem_arlock,
  output [3:0]  io_mem_arcache,
  output [3:0]  io_mem_arqos,
  output        io_mem_rready,
  input         io_mem_rvalid,
  input  [1:0]  io_mem_rresp,
  input  [63:0] io_mem_rdata,
  input         io_mem_rlast,
  input         io_mem_rid,
  input         io_mem_ruser,
  input         io_mmio_awready,
  output        io_mmio_awvalid,
  output [31:0] io_mmio_awaddr,
  output [2:0]  io_mmio_awprot,
  output        io_mmio_awid,
  output        io_mmio_awuser,
  output [7:0]  io_mmio_awlen,
  output [2:0]  io_mmio_awsize,
  output [1:0]  io_mmio_awburst,
  output        io_mmio_awlock,
  output [3:0]  io_mmio_awcache,
  output [3:0]  io_mmio_awqos,
  input         io_mmio_wready,
  output        io_mmio_wvalid,
  output [63:0] io_mmio_wdata,
  output [7:0]  io_mmio_wstrb,
  output        io_mmio_wlast,
  output        io_mmio_bready,
  input         io_mmio_bvalid,
  input  [1:0]  io_mmio_bresp,
  input         io_mmio_bid,
  input         io_mmio_buser,
  input         io_mmio_arready,
  output        io_mmio_arvalid,
  output [31:0] io_mmio_araddr,
  output [2:0]  io_mmio_arprot,
  output        io_mmio_arid,
  output        io_mmio_aruser,
  output [7:0]  io_mmio_arlen,
  output [2:0]  io_mmio_arsize,
  output [1:0]  io_mmio_arburst,
  output        io_mmio_arlock,
  output [3:0]  io_mmio_arcache,
  output [3:0]  io_mmio_arqos,
  output        io_mmio_rready,
  input         io_mmio_rvalid,
  input  [1:0]  io_mmio_rresp,
  input  [63:0] io_mmio_rdata,
  input         io_mmio_rlast,
  input         io_mmio_rid,
  input         io_mmio_ruser,
  output        io_frontend_awready,
  input         io_frontend_awvalid,
  input  [31:0] io_frontend_awaddr,
  input  [2:0]  io_frontend_awprot,
  input         io_frontend_awid,
  input         io_frontend_awuser,
  input  [7:0]  io_frontend_awlen,
  input  [2:0]  io_frontend_awsize,
  input  [1:0]  io_frontend_awburst,
  input         io_frontend_awlock,
  input  [3:0]  io_frontend_awcache,
  input  [3:0]  io_frontend_awqos,
  output        io_frontend_wready,
  input         io_frontend_wvalid,
  input  [63:0] io_frontend_wdata,
  input  [7:0]  io_frontend_wstrb,
  input         io_frontend_wlast,
  input         io_frontend_bready,
  output        io_frontend_bvalid,
  output [1:0]  io_frontend_bresp,
  output        io_frontend_bid,
  output        io_frontend_buser,
  output        io_frontend_arready,
  input         io_frontend_arvalid,
  input  [31:0] io_frontend_araddr,
  input  [2:0]  io_frontend_arprot,
  input         io_frontend_arid,
  input         io_frontend_aruser,
  input  [7:0]  io_frontend_arlen,
  input  [2:0]  io_frontend_arsize,
  input  [1:0]  io_frontend_arburst,
  input         io_frontend_arlock,
  input  [3:0]  io_frontend_arcache,
  input  [3:0]  io_frontend_arqos,
  input         io_frontend_rready,
  output        io_frontend_rvalid,
  output [1:0]  io_frontend_rresp,
  output [63:0] io_frontend_rdata,
  output        io_frontend_rlast,
  output        io_frontend_rid,
  output        io_frontend_ruser,
  input  [2:0]  io_meip,
  output [38:0] io_ila_WBUpc,
  output        io_ila_WBUvalid,
  output        io_ila_WBUrfWen,
  output [4:0]  io_ila_WBUrfDest,
  output [63:0] io_ila_WBUrfData,
  output [63:0] io_ila_InstrCnt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  nutcore_clock; // @[NutShell.scala 53:23]
  wire  nutcore_reset; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_coh_req_bits_addr; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_mmio_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_frontend_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_frontend_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_frontend_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_perfCnts_2; // @[NutShell.scala 53:23]
  wire [38:0] nutcore_io_in_0_bits_decode_cf_pc; // @[NutShell.scala 53:23]
  wire [4:0] nutcore_io_wb_rfDest_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_wb_rfWen_0; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_wb_WriteData_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[NutShell.scala 53:23]
  wire  nutcore_io_in_0_valid_0; // @[NutShell.scala 53:23]
  wire  cohMg_clock; // @[NutShell.scala 54:21]
  wire  cohMg_reset; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_coh_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  xbar_clock; // @[NutShell.scala 55:20]
  wire  xbar_reset; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_in_0_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_0_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  axi2sb_clock; // @[NutShell.scala 61:22]
  wire  axi2sb_reset; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_awready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_awvalid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_awaddr; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_awid; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_awlen; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_awsize; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wvalid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_wdata; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_wstrb; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wlast; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_bready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_bvalid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_arready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_arvalid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_araddr; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_arid; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_arlen; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_arsize; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rvalid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_rdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rlast; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_rid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_valid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_out_req_bits_addr; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_out_req_bits_size; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_valid; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_resp_bits_cmd; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_resp_bits_rdata; // @[NutShell.scala 61:22]
  wire  Prefetcher_clock; // @[NutShell.scala 73:30]
  wire  Prefetcher_reset; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_in_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_in_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_in_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_in_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_in_bits_wdata; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_out_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_out_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_out_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_out_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_out_bits_wdata; // @[NutShell.scala 73:30]
  wire  Cache_clock; // @[Cache.scala 674:35]
  wire  Cache_reset; // @[Cache.scala 674:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 674:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 674:35]
  wire [2:0] Cache_io_in_req_bits_size; // @[Cache.scala 674:35]
  wire [3:0] Cache_io_in_req_bits_cmd; // @[Cache.scala 674:35]
  wire [7:0] Cache_io_in_req_bits_wmask; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_in_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 674:35]
  wire [3:0] Cache_io_in_resp_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 674:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 674:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 674:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 674:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 674:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 674:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 674:35]
  wire  memAddrMap_io_in_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  SimpleBus2AXI4Converter_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awuser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aruser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_in_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_2_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  SimpleBus2AXI4Converter_1_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_in_req_bits_size; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_awprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awuser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_1_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_awcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_awqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_arprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aruser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_1_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_arcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_arqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  clint_clock; // @[NutShell.scala 113:21]
  wire  clint_reset; // @[NutShell.scala 113:21]
  wire  clint_io__in_awready; // @[NutShell.scala 113:21]
  wire  clint_io__in_awvalid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_awaddr; // @[NutShell.scala 113:21]
  wire  clint_io__in_wready; // @[NutShell.scala 113:21]
  wire  clint_io__in_wvalid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_wdata; // @[NutShell.scala 113:21]
  wire [7:0] clint_io__in_wstrb; // @[NutShell.scala 113:21]
  wire  clint_io__in_bready; // @[NutShell.scala 113:21]
  wire  clint_io__in_bvalid; // @[NutShell.scala 113:21]
  wire  clint_io__in_arready; // @[NutShell.scala 113:21]
  wire  clint_io__in_arvalid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_araddr; // @[NutShell.scala 113:21]
  wire  clint_io__in_rready; // @[NutShell.scala 113:21]
  wire  clint_io__in_rvalid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_rdata; // @[NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[NutShell.scala 113:21]
  wire  SimpleBus2AXI4Converter_2_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_2_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  plic_clock; // @[NutShell.scala 120:20]
  wire  plic_reset; // @[NutShell.scala 120:20]
  wire  plic_io__in_awready; // @[NutShell.scala 120:20]
  wire  plic_io__in_awvalid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_awaddr; // @[NutShell.scala 120:20]
  wire  plic_io__in_wready; // @[NutShell.scala 120:20]
  wire  plic_io__in_wvalid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_wdata; // @[NutShell.scala 120:20]
  wire [7:0] plic_io__in_wstrb; // @[NutShell.scala 120:20]
  wire  plic_io__in_bready; // @[NutShell.scala 120:20]
  wire  plic_io__in_bvalid; // @[NutShell.scala 120:20]
  wire  plic_io__in_arready; // @[NutShell.scala 120:20]
  wire  plic_io__in_arvalid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_araddr; // @[NutShell.scala 120:20]
  wire  plic_io__in_rready; // @[NutShell.scala 120:20]
  wire  plic_io__in_rvalid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_rdata; // @[NutShell.scala 120:20]
  wire [2:0] plic_io__extra_intrVec; // @[NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[NutShell.scala 120:20]
  wire  SimpleBus2AXI4Converter_3_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_3_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_rdata; // @[ToAXI4.scala 204:24]
  reg [2:0] REG; // @[NutShell.scala 122:47]
  reg [2:0] REG_1; // @[NutShell.scala 122:39]
  wire  ilaWBUvalid = nutcore_io_in_0_valid_0;
  wire  ilaWBUrfWen = nutcore_io_wb_rfWen_0;
  wire [4:0] ilaWBUrfDest = nutcore_io_wb_rfDest_0;
  wire [38:0] ilaWBUpc = nutcore_io_in_0_bits_decode_cf_pc;
  wire [63:0] _WIRE_6 = {{25'd0}, ilaWBUpc};
  wire [63:0] _WIRE_7 = {{63'd0}, ilaWBUvalid};
  wire [63:0] _WIRE_8 = {{63'd0}, ilaWBUrfWen};
  wire [63:0] _WIRE_9 = {{59'd0}, ilaWBUrfDest};
  NutCore nutcore ( // @[NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_req_bits_cmd(nutcore_io_imem_mem_req_bits_cmd),
    .io_imem_mem_req_bits_wdata(nutcore_io_imem_mem_req_bits_wdata),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_cmd(nutcore_io_imem_mem_resp_bits_cmd),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_dmem_coh_req_ready(nutcore_io_dmem_coh_req_ready),
    .io_dmem_coh_req_valid(nutcore_io_dmem_coh_req_valid),
    .io_dmem_coh_req_bits_addr(nutcore_io_dmem_coh_req_bits_addr),
    .io_dmem_coh_req_bits_wdata(nutcore_io_dmem_coh_req_bits_wdata),
    .io_dmem_coh_resp_valid(nutcore_io_dmem_coh_resp_valid),
    .io_dmem_coh_resp_bits_cmd(nutcore_io_dmem_coh_resp_bits_cmd),
    .io_dmem_coh_resp_bits_rdata(nutcore_io_dmem_coh_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(nutcore_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_frontend_req_valid(nutcore_io_frontend_req_valid),
    .io_frontend_req_bits_addr(nutcore_io_frontend_req_bits_addr),
    .io_frontend_req_bits_size(nutcore_io_frontend_req_bits_size),
    .io_frontend_req_bits_cmd(nutcore_io_frontend_req_bits_cmd),
    .io_frontend_req_bits_wmask(nutcore_io_frontend_req_bits_wmask),
    .io_frontend_req_bits_wdata(nutcore_io_frontend_req_bits_wdata),
    .io_frontend_resp_ready(nutcore_io_frontend_resp_ready),
    .io_frontend_resp_valid(nutcore_io_frontend_resp_valid),
    .io_frontend_resp_bits_cmd(nutcore_io_frontend_resp_bits_cmd),
    .io_frontend_resp_bits_rdata(nutcore_io_frontend_resp_bits_rdata),
    .perfCnts_2(nutcore_perfCnts_2),
    .io_in_0_bits_decode_cf_pc(nutcore_io_in_0_bits_decode_cf_pc),
    .io_wb_rfDest_0(nutcore_io_wb_rfDest_0),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .io_wb_rfWen_0(nutcore_io_wb_rfWen_0),
    .io_wb_WriteData_0(nutcore_io_wb_WriteData_0),
    .io_extra_msip(nutcore_io_extra_msip),
    .io_in_0_valid_0(nutcore_io_in_0_valid_0)
  );
  CoherenceManager cohMg ( // @[NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_req_bits_cmd(cohMg_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(cohMg_io_in_req_bits_wdata),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(cohMg_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(cohMg_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(cohMg_io_out_coh_req_ready),
    .io_out_coh_req_valid(cohMg_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(cohMg_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(cohMg_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_ready(cohMg_io_out_coh_resp_ready),
    .io_out_coh_resp_valid(cohMg_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(cohMg_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(cohMg_io_out_coh_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1 xbar ( // @[NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(xbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(xbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(xbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(xbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_in_awready(axi2sb_io_in_awready),
    .io_in_awvalid(axi2sb_io_in_awvalid),
    .io_in_awaddr(axi2sb_io_in_awaddr),
    .io_in_awid(axi2sb_io_in_awid),
    .io_in_awlen(axi2sb_io_in_awlen),
    .io_in_awsize(axi2sb_io_in_awsize),
    .io_in_wready(axi2sb_io_in_wready),
    .io_in_wvalid(axi2sb_io_in_wvalid),
    .io_in_wdata(axi2sb_io_in_wdata),
    .io_in_wstrb(axi2sb_io_in_wstrb),
    .io_in_wlast(axi2sb_io_in_wlast),
    .io_in_bready(axi2sb_io_in_bready),
    .io_in_bvalid(axi2sb_io_in_bvalid),
    .io_in_arready(axi2sb_io_in_arready),
    .io_in_arvalid(axi2sb_io_in_arvalid),
    .io_in_araddr(axi2sb_io_in_araddr),
    .io_in_arid(axi2sb_io_in_arid),
    .io_in_arlen(axi2sb_io_in_arlen),
    .io_in_arsize(axi2sb_io_in_arsize),
    .io_in_rready(axi2sb_io_in_rready),
    .io_in_rvalid(axi2sb_io_in_rvalid),
    .io_in_rdata(axi2sb_io_in_rdata),
    .io_in_rlast(axi2sb_io_in_rlast),
    .io_in_rid(axi2sb_io_in_rid),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid),
    .io_out_req_bits_addr(axi2sb_io_out_req_bits_addr),
    .io_out_req_bits_size(axi2sb_io_out_req_bits_size),
    .io_out_req_bits_cmd(axi2sb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(axi2sb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(axi2sb_io_out_req_bits_wdata),
    .io_out_resp_ready(axi2sb_io_out_resp_ready),
    .io_out_resp_valid(axi2sb_io_out_resp_valid),
    .io_out_resp_bits_cmd(axi2sb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(axi2sb_io_out_resp_bits_rdata)
  );
  Prefetcher Prefetcher ( // @[NutShell.scala 73:30]
    .clock(Prefetcher_clock),
    .reset(Prefetcher_reset),
    .io_in_ready(Prefetcher_io_in_ready),
    .io_in_valid(Prefetcher_io_in_valid),
    .io_in_bits_addr(Prefetcher_io_in_bits_addr),
    .io_in_bits_size(Prefetcher_io_in_bits_size),
    .io_in_bits_cmd(Prefetcher_io_in_bits_cmd),
    .io_in_bits_wmask(Prefetcher_io_in_bits_wmask),
    .io_in_bits_wdata(Prefetcher_io_in_bits_wdata),
    .io_out_ready(Prefetcher_io_out_ready),
    .io_out_valid(Prefetcher_io_out_valid),
    .io_out_bits_addr(Prefetcher_io_out_bits_addr),
    .io_out_bits_size(Prefetcher_io_out_bits_size),
    .io_out_bits_cmd(Prefetcher_io_out_bits_cmd),
    .io_out_bits_wmask(Prefetcher_io_out_bits_wmask),
    .io_out_bits_wdata(Prefetcher_io_out_bits_wdata)
  );
  Cache_2 Cache ( // @[Cache.scala 674:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_io_in_req_bits_wdata),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata)
  );
  SimpleBusAddressMapper memAddrMap ( // @[NutShell.scala 93:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter SimpleBus2AXI4Converter ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_clock),
    .reset(SimpleBus2AXI4Converter_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_io_in_req_bits_wdata),
    .io_in_resp_valid(SimpleBus2AXI4Converter_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_io_out_awaddr),
    .io_out_awprot(SimpleBus2AXI4Converter_io_out_awprot),
    .io_out_awid(SimpleBus2AXI4Converter_io_out_awid),
    .io_out_awuser(SimpleBus2AXI4Converter_io_out_awuser),
    .io_out_awlen(SimpleBus2AXI4Converter_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_io_out_awburst),
    .io_out_awlock(SimpleBus2AXI4Converter_io_out_awlock),
    .io_out_awcache(SimpleBus2AXI4Converter_io_out_awcache),
    .io_out_awqos(SimpleBus2AXI4Converter_io_out_awqos),
    .io_out_wready(SimpleBus2AXI4Converter_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_io_out_wdata),
    .io_out_wlast(SimpleBus2AXI4Converter_io_out_wlast),
    .io_out_bvalid(SimpleBus2AXI4Converter_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_io_out_araddr),
    .io_out_arprot(SimpleBus2AXI4Converter_io_out_arprot),
    .io_out_arid(SimpleBus2AXI4Converter_io_out_arid),
    .io_out_aruser(SimpleBus2AXI4Converter_io_out_aruser),
    .io_out_arlen(SimpleBus2AXI4Converter_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_io_out_arburst),
    .io_out_arlock(SimpleBus2AXI4Converter_io_out_arlock),
    .io_out_arcache(SimpleBus2AXI4Converter_io_out_arcache),
    .io_out_arqos(SimpleBus2AXI4Converter_io_out_arqos),
    .io_out_rvalid(SimpleBus2AXI4Converter_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_io_out_rlast)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_size(mmioXbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_size(mmioXbar_io_out_2_req_bits_size),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_cmd(mmioXbar_io_out_2_resp_bits_cmd),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_1 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_1_clock),
    .reset(SimpleBus2AXI4Converter_1_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_1_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_1_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_1_io_in_req_bits_addr),
    .io_in_req_bits_size(SimpleBus2AXI4Converter_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_1_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_1_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_1_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_1_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_1_io_out_awaddr),
    .io_out_awprot(SimpleBus2AXI4Converter_1_io_out_awprot),
    .io_out_awid(SimpleBus2AXI4Converter_1_io_out_awid),
    .io_out_awuser(SimpleBus2AXI4Converter_1_io_out_awuser),
    .io_out_awlen(SimpleBus2AXI4Converter_1_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_1_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_1_io_out_awburst),
    .io_out_awlock(SimpleBus2AXI4Converter_1_io_out_awlock),
    .io_out_awcache(SimpleBus2AXI4Converter_1_io_out_awcache),
    .io_out_awqos(SimpleBus2AXI4Converter_1_io_out_awqos),
    .io_out_wready(SimpleBus2AXI4Converter_1_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_1_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_1_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_1_io_out_wstrb),
    .io_out_wlast(SimpleBus2AXI4Converter_1_io_out_wlast),
    .io_out_bready(SimpleBus2AXI4Converter_1_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_1_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_1_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_1_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_1_io_out_araddr),
    .io_out_arprot(SimpleBus2AXI4Converter_1_io_out_arprot),
    .io_out_arid(SimpleBus2AXI4Converter_1_io_out_arid),
    .io_out_aruser(SimpleBus2AXI4Converter_1_io_out_aruser),
    .io_out_arlen(SimpleBus2AXI4Converter_1_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_1_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_1_io_out_arburst),
    .io_out_arlock(SimpleBus2AXI4Converter_1_io_out_arlock),
    .io_out_arcache(SimpleBus2AXI4Converter_1_io_out_arcache),
    .io_out_arqos(SimpleBus2AXI4Converter_1_io_out_arqos),
    .io_out_rready(SimpleBus2AXI4Converter_1_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_1_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_1_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_1_io_out_rlast)
  );
  AXI4CLINT clint ( // @[NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_awready(clint_io__in_awready),
    .io__in_awvalid(clint_io__in_awvalid),
    .io__in_awaddr(clint_io__in_awaddr),
    .io__in_wready(clint_io__in_wready),
    .io__in_wvalid(clint_io__in_wvalid),
    .io__in_wdata(clint_io__in_wdata),
    .io__in_wstrb(clint_io__in_wstrb),
    .io__in_bready(clint_io__in_bready),
    .io__in_bvalid(clint_io__in_bvalid),
    .io__in_arready(clint_io__in_arready),
    .io__in_arvalid(clint_io__in_arvalid),
    .io__in_araddr(clint_io__in_araddr),
    .io__in_rready(clint_io__in_rready),
    .io__in_rvalid(clint_io__in_rvalid),
    .io__in_rdata(clint_io__in_rdata),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_2 SimpleBus2AXI4Converter_2 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_2_clock),
    .reset(SimpleBus2AXI4Converter_2_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_2_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_2_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_2_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_2_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_2_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_2_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_2_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_2_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_2_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_2_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_2_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_2_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_2_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_2_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_2_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_2_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_2_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_2_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_2_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_2_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_2_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_2_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_2_io_out_rdata)
  );
  AXI4PLIC plic ( // @[NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_awready(plic_io__in_awready),
    .io__in_awvalid(plic_io__in_awvalid),
    .io__in_awaddr(plic_io__in_awaddr),
    .io__in_wready(plic_io__in_wready),
    .io__in_wvalid(plic_io__in_wvalid),
    .io__in_wdata(plic_io__in_wdata),
    .io__in_wstrb(plic_io__in_wstrb),
    .io__in_bready(plic_io__in_bready),
    .io__in_bvalid(plic_io__in_bvalid),
    .io__in_arready(plic_io__in_arready),
    .io__in_arvalid(plic_io__in_arvalid),
    .io__in_araddr(plic_io__in_araddr),
    .io__in_rready(plic_io__in_rready),
    .io__in_rvalid(plic_io__in_rvalid),
    .io__in_rdata(plic_io__in_rdata),
    .io__extra_intrVec(plic_io__extra_intrVec),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_2 SimpleBus2AXI4Converter_3 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_3_clock),
    .reset(SimpleBus2AXI4Converter_3_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_3_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_3_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_3_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_3_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_3_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_3_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_3_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_3_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_3_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_3_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_3_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_3_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_3_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_3_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_3_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_3_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_3_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_3_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_3_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_3_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_3_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_3_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_3_io_out_rdata)
  );
  assign io_mem_awvalid = SimpleBus2AXI4Converter_io_out_awvalid; // @[NutShell.scala 95:10]
  assign io_mem_awaddr = SimpleBus2AXI4Converter_io_out_awaddr; // @[NutShell.scala 95:10]
  assign io_mem_awprot = SimpleBus2AXI4Converter_io_out_awprot; // @[NutShell.scala 95:10]
  assign io_mem_awid = SimpleBus2AXI4Converter_io_out_awid; // @[NutShell.scala 95:10]
  assign io_mem_awuser = SimpleBus2AXI4Converter_io_out_awuser; // @[NutShell.scala 95:10]
  assign io_mem_awlen = SimpleBus2AXI4Converter_io_out_awlen; // @[NutShell.scala 95:10]
  assign io_mem_awsize = SimpleBus2AXI4Converter_io_out_awsize; // @[NutShell.scala 95:10]
  assign io_mem_awburst = SimpleBus2AXI4Converter_io_out_awburst; // @[NutShell.scala 95:10]
  assign io_mem_awlock = SimpleBus2AXI4Converter_io_out_awlock; // @[NutShell.scala 95:10]
  assign io_mem_awcache = SimpleBus2AXI4Converter_io_out_awcache; // @[NutShell.scala 95:10]
  assign io_mem_awqos = SimpleBus2AXI4Converter_io_out_awqos; // @[NutShell.scala 95:10]
  assign io_mem_wvalid = SimpleBus2AXI4Converter_io_out_wvalid; // @[NutShell.scala 95:10]
  assign io_mem_wdata = SimpleBus2AXI4Converter_io_out_wdata; // @[NutShell.scala 95:10]
  assign io_mem_wstrb = 8'hff; // @[NutShell.scala 95:10]
  assign io_mem_wlast = SimpleBus2AXI4Converter_io_out_wlast; // @[NutShell.scala 95:10]
  assign io_mem_bready = 1'h1; // @[NutShell.scala 95:10]
  assign io_mem_arvalid = SimpleBus2AXI4Converter_io_out_arvalid; // @[NutShell.scala 95:10]
  assign io_mem_araddr = SimpleBus2AXI4Converter_io_out_araddr; // @[NutShell.scala 95:10]
  assign io_mem_arprot = 3'h1; // @[NutShell.scala 95:10]
  assign io_mem_arid = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_aruser = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_arlen = SimpleBus2AXI4Converter_io_out_arlen; // @[NutShell.scala 95:10]
  assign io_mem_arsize = 3'h3; // @[NutShell.scala 95:10]
  assign io_mem_arburst = 2'h2; // @[NutShell.scala 95:10]
  assign io_mem_arlock = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_arcache = 4'h0; // @[NutShell.scala 95:10]
  assign io_mem_arqos = 4'h0; // @[NutShell.scala 95:10]
  assign io_mem_rready = 1'h1; // @[NutShell.scala 95:10]
  assign io_mmio_awvalid = SimpleBus2AXI4Converter_1_io_out_awvalid; // @[NutShell.scala 110:33]
  assign io_mmio_awaddr = SimpleBus2AXI4Converter_1_io_out_awaddr; // @[NutShell.scala 110:33]
  assign io_mmio_awprot = SimpleBus2AXI4Converter_1_io_out_awprot; // @[NutShell.scala 110:33]
  assign io_mmio_awid = SimpleBus2AXI4Converter_1_io_out_awid; // @[NutShell.scala 110:33]
  assign io_mmio_awuser = SimpleBus2AXI4Converter_1_io_out_awuser; // @[NutShell.scala 110:33]
  assign io_mmio_awlen = SimpleBus2AXI4Converter_1_io_out_awlen; // @[NutShell.scala 110:33]
  assign io_mmio_awsize = SimpleBus2AXI4Converter_1_io_out_awsize; // @[NutShell.scala 110:33]
  assign io_mmio_awburst = SimpleBus2AXI4Converter_1_io_out_awburst; // @[NutShell.scala 110:33]
  assign io_mmio_awlock = SimpleBus2AXI4Converter_1_io_out_awlock; // @[NutShell.scala 110:33]
  assign io_mmio_awcache = SimpleBus2AXI4Converter_1_io_out_awcache; // @[NutShell.scala 110:33]
  assign io_mmio_awqos = SimpleBus2AXI4Converter_1_io_out_awqos; // @[NutShell.scala 110:33]
  assign io_mmio_wvalid = SimpleBus2AXI4Converter_1_io_out_wvalid; // @[NutShell.scala 110:33]
  assign io_mmio_wdata = SimpleBus2AXI4Converter_1_io_out_wdata; // @[NutShell.scala 110:33]
  assign io_mmio_wstrb = SimpleBus2AXI4Converter_1_io_out_wstrb; // @[NutShell.scala 110:33]
  assign io_mmio_wlast = SimpleBus2AXI4Converter_1_io_out_wlast; // @[NutShell.scala 110:33]
  assign io_mmio_bready = SimpleBus2AXI4Converter_1_io_out_bready; // @[NutShell.scala 110:33]
  assign io_mmio_arvalid = SimpleBus2AXI4Converter_1_io_out_arvalid; // @[NutShell.scala 110:33]
  assign io_mmio_araddr = SimpleBus2AXI4Converter_1_io_out_araddr; // @[NutShell.scala 110:33]
  assign io_mmio_arprot = 3'h1; // @[NutShell.scala 110:33]
  assign io_mmio_arid = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_aruser = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arlen = SimpleBus2AXI4Converter_1_io_out_arlen; // @[NutShell.scala 110:33]
  assign io_mmio_arsize = SimpleBus2AXI4Converter_1_io_out_arsize; // @[NutShell.scala 110:33]
  assign io_mmio_arburst = 2'h1; // @[NutShell.scala 110:33]
  assign io_mmio_arlock = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arcache = 4'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arqos = 4'h0; // @[NutShell.scala 110:33]
  assign io_mmio_rready = SimpleBus2AXI4Converter_1_io_out_rready; // @[NutShell.scala 110:33]
  assign io_frontend_awready = axi2sb_io_in_awready; // @[NutShell.scala 62:16]
  assign io_frontend_wready = axi2sb_io_in_wready; // @[NutShell.scala 62:16]
  assign io_frontend_bvalid = axi2sb_io_in_bvalid; // @[NutShell.scala 62:16]
  assign io_frontend_bresp = 2'h0; // @[NutShell.scala 62:16]
  assign io_frontend_bid = 1'h0; // @[NutShell.scala 62:16]
  assign io_frontend_buser = 1'h0; // @[NutShell.scala 62:16]
  assign io_frontend_arready = axi2sb_io_in_arready; // @[NutShell.scala 62:16]
  assign io_frontend_rvalid = axi2sb_io_in_rvalid; // @[NutShell.scala 62:16]
  assign io_frontend_rresp = 2'h0; // @[NutShell.scala 62:16]
  assign io_frontend_rdata = axi2sb_io_in_rdata; // @[NutShell.scala 62:16]
  assign io_frontend_rlast = axi2sb_io_in_rlast; // @[NutShell.scala 62:16]
  assign io_frontend_rid = axi2sb_io_in_rid[0]; // @[NutShell.scala 62:16]
  assign io_frontend_ruser = 1'h0; // @[NutShell.scala 62:16]
  assign io_ila_WBUpc = _WIRE_6[38:0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUvalid = _WIRE_7[0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfWen = _WIRE_8[0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfDest = _WIRE_9[4:0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfData = nutcore_io_wb_WriteData_0; // @[NutShell.scala 132:12]
  assign io_ila_InstrCnt = nutcore_perfCnts_2; // @[NutShell.scala 132:12]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_cmd = cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_coh_req_valid = cohMg_io_out_coh_req_valid; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_addr = cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_wdata = cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 57:23]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 107:18]
  assign nutcore_io_frontend_req_valid = axi2sb_io_out_req_valid; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_addr = axi2sb_io_out_req_bits_addr; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_size = axi2sb_io_out_req_bits_size; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_cmd = axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wmask = axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wdata = axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_resp_ready = axi2sb_io_out_resp_ready; // @[NutShell.scala 63:23]
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_cmd = nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_wdata = nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 58:17]
  assign cohMg_io_out_coh_req_ready = nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_valid = nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_cmd = nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_rdata = nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 57:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_size = 3'h3; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_cmd = cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wmask = 8'hff; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wdata = cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = 3'h3; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = 8'hff; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 59:17]
  assign xbar_io_out_req_ready = Prefetcher_io_in_ready; // @[NutShell.scala 75:24]
  assign xbar_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 680:17 NutShell.scala 74:27]
  assign xbar_io_out_resp_bits_cmd = Cache_io_in_resp_bits_cmd; // @[Cache.scala 680:17 NutShell.scala 74:27]
  assign xbar_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 680:17 NutShell.scala 74:27]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_in_awvalid = io_frontend_awvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awaddr = io_frontend_awaddr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awid = {{17'd0}, io_frontend_awid}; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awlen = io_frontend_awlen; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awsize = io_frontend_awsize; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wvalid = io_frontend_wvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wdata = io_frontend_wdata; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wstrb = io_frontend_wstrb; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wlast = io_frontend_wlast; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_bready = io_frontend_bready; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arvalid = io_frontend_arvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_araddr = io_frontend_araddr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arid = {{17'd0}, io_frontend_arid}; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arlen = io_frontend_arlen; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arsize = io_frontend_arsize; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_rready = io_frontend_rready; // @[NutShell.scala 62:16]
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_valid = nutcore_io_frontend_resp_valid; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_cmd = nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_rdata = nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 63:23]
  assign Prefetcher_clock = clock;
  assign Prefetcher_reset = reset;
  assign Prefetcher_io_in_valid = xbar_io_out_req_valid; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_addr = xbar_io_out_req_bits_addr; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_size = xbar_io_out_req_bits_size; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_cmd = xbar_io_out_req_bits_cmd; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wmask = xbar_io_out_req_bits_wmask; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wdata = xbar_io_out_req_bits_wdata; // @[NutShell.scala 75:24]
  assign Prefetcher_io_out_ready = Cache_io_in_req_ready; // @[Cache.scala 680:17 NutShell.scala 74:27]
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = Prefetcher_io_out_valid; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_addr = Prefetcher_io_out_bits_addr; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_size = Prefetcher_io_out_bits_size; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_cmd = Prefetcher_io_out_bits_cmd; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_wmask = Prefetcher_io_out_bits_wmask; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_wdata = Prefetcher_io_out_bits_wdata; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_out_mem_req_ready = memAddrMap_io_in_req_ready; // @[NutShell.scala 71:26 94:20]
  assign Cache_io_out_mem_resp_valid = memAddrMap_io_in_resp_valid; // @[NutShell.scala 71:26 94:20]
  assign Cache_io_out_mem_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 71:26 94:20]
  assign Cache_io_out_mem_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 71:26 94:20]
  assign memAddrMap_io_in_req_valid = Cache_io_out_mem_req_valid; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_out_req_ready = SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_clock = clock;
  assign SimpleBus2AXI4Converter_reset = reset;
  assign SimpleBus2AXI4Converter_io_in_req_valid = memAddrMap_io_out_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_out_awready = io_mem_awready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_wready = io_mem_wready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_bvalid = io_mem_bvalid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_arready = io_mem_arready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rvalid = io_mem_rvalid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rdata = io_mem_rdata; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rlast = io_mem_rlast; // @[NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_size = nutcore_io_mmio_req_bits_size; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_valid = SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_bits_cmd = SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_clock = clock;
  assign SimpleBus2AXI4Converter_1_reset = reset;
  assign SimpleBus2AXI4Converter_1_io_in_req_valid = mmioXbar_io_out_2_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_size = mmioXbar_io_out_2_req_bits_size; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_resp_ready = mmioXbar_io_out_2_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_out_awready = io_mmio_awready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_wready = io_mmio_wready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_bvalid = io_mmio_bvalid; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_arready = io_mmio_arready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rvalid = io_mmio_rvalid; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rdata = io_mmio_rdata; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rlast = io_mmio_rlast; // @[NutShell.scala 110:33]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_awvalid = SimpleBus2AXI4Converter_2_io_out_awvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_awaddr = SimpleBus2AXI4Converter_2_io_out_awaddr; // @[NutShell.scala 114:15]
  assign clint_io__in_wvalid = SimpleBus2AXI4Converter_2_io_out_wvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_wdata = SimpleBus2AXI4Converter_2_io_out_wdata; // @[NutShell.scala 114:15]
  assign clint_io__in_wstrb = SimpleBus2AXI4Converter_2_io_out_wstrb; // @[NutShell.scala 114:15]
  assign clint_io__in_bready = SimpleBus2AXI4Converter_2_io_out_bready; // @[NutShell.scala 114:15]
  assign clint_io__in_arvalid = SimpleBus2AXI4Converter_2_io_out_arvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_araddr = SimpleBus2AXI4Converter_2_io_out_araddr; // @[NutShell.scala 114:15]
  assign clint_io__in_rready = SimpleBus2AXI4Converter_2_io_out_rready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_clock = clock;
  assign SimpleBus2AXI4Converter_2_reset = reset;
  assign SimpleBus2AXI4Converter_2_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_out_awready = clint_io__in_awready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_wready = clint_io__in_wready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_bvalid = clint_io__in_bvalid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_arready = clint_io__in_arready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_rvalid = clint_io__in_rvalid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_rdata = clint_io__in_rdata; // @[NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_awvalid = SimpleBus2AXI4Converter_3_io_out_awvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_awaddr = SimpleBus2AXI4Converter_3_io_out_awaddr; // @[NutShell.scala 121:14]
  assign plic_io__in_wvalid = SimpleBus2AXI4Converter_3_io_out_wvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_wdata = SimpleBus2AXI4Converter_3_io_out_wdata; // @[NutShell.scala 121:14]
  assign plic_io__in_wstrb = SimpleBus2AXI4Converter_3_io_out_wstrb; // @[NutShell.scala 121:14]
  assign plic_io__in_bready = SimpleBus2AXI4Converter_3_io_out_bready; // @[NutShell.scala 121:14]
  assign plic_io__in_arvalid = SimpleBus2AXI4Converter_3_io_out_arvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_araddr = SimpleBus2AXI4Converter_3_io_out_araddr; // @[NutShell.scala 121:14]
  assign plic_io__in_rready = SimpleBus2AXI4Converter_3_io_out_rready; // @[NutShell.scala 121:14]
  assign plic_io__extra_intrVec = REG_1; // @[NutShell.scala 122:29]
  assign SimpleBus2AXI4Converter_3_clock = clock;
  assign SimpleBus2AXI4Converter_3_reset = reset;
  assign SimpleBus2AXI4Converter_3_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_out_awready = plic_io__in_awready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_wready = plic_io__in_wready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_bvalid = plic_io__in_bvalid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_arready = plic_io__in_arready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_rvalid = plic_io__in_rvalid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_rdata = plic_io__in_rdata; // @[NutShell.scala 121:14]
  always @(posedge clock) begin
    REG <= io_meip; // @[NutShell.scala 122:47]
    REG_1 <= REG; // @[NutShell.scala 122:39]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  output        io_in_wready,
  input         io_in_wvalid,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  _T_24 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_25 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_25 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_25 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  wire  _T_73 = 4'h0 == io_in_araddr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_74 = 4'h4 == io_in_araddr[3:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_75 = _T_73 ? 32'h190012c : 32'h0; // @[Mux.scala 27:72]
  wire  _T_76 = _T_74 & _T_38; // @[Mux.scala 27:72]
  wire [31:0] _GEN_8 = {{31'd0}, _T_76}; // @[Mux.scala 27:72]
  wire [31:0] _T_77 = _T_75 | _GEN_8; // @[Mux.scala 27:72]
  assign io_in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io_in_wready = io_in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io_in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io_in_arready = io_in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io_in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io_in_rdata = {{32'd0}, _T_77}; // @[RegMap.scala 30:11]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] MEM_0 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_0_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_0_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_0_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_0_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_0_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_0_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_0_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_1 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_1_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_1_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_1_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_1_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_1_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_1_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_1_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_2 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_2_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_2_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_2_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_2_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_2_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_2_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_2_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_3 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_3_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_3_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_3_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_3_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_3_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_3_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_3_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_4 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_4_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_4_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_4_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_4_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_4_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_4_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_4_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_5 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_5_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_5_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_5_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_5_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_5_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_5_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_5_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_6 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_6_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_6_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_6_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_6_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_6_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_6_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_6_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_7 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_7_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_7_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_7_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_7_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_7_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_7_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_7_MPORT_en; // @[AXI4RAM.scala 63:18]
  wire  _T_24 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_rvalid ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = io_in_rvalid ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  wire [31:0] _T_45 = io_in_awaddr & 32'h7ffff; // @[AXI4RAM.scala 45:33]
  wire [29:0] _T_47 = {{1'd0}, _T_45[31:3]}; // @[AXI4RAM.scala 48:27]
  wire [28:0] wIdx = _T_47[28:0]; // @[AXI4RAM.scala 48:27]
  wire [31:0] _T_48 = io_in_araddr & 32'h7ffff; // @[AXI4RAM.scala 45:33]
  wire [29:0] _T_50 = {{1'd0}, _T_48[31:3]}; // @[AXI4RAM.scala 49:27]
  wire [28:0] rIdx = _T_50[28:0]; // @[AXI4RAM.scala 49:27]
  wire  _T_52 = wIdx < 29'hea60; // @[AXI4RAM.scala 46:32]
  wire [63:0] rdata = {MEM_7_MPORT_1_data,MEM_6_MPORT_1_data,MEM_5_MPORT_1_data,MEM_4_MPORT_1_data,MEM_3_MPORT_1_data,
    MEM_2_MPORT_1_data,MEM_1_MPORT_1_data,MEM_0_MPORT_1_data}; // @[Cat.scala 30:58]
  reg [63:0] r; // @[Reg.scala 15:16]
  assign MEM_0_MPORT_1_en = 1'h1;
  assign MEM_0_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_0_MPORT_1_data = MEM_0[MEM_0_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_0_MPORT_1_data = MEM_0_MPORT_1_addr >= 16'hea60 ? _RAND_1[7:0] : MEM_0[MEM_0_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_0_MPORT_data = io_in_wdata[7:0];
  assign MEM_0_MPORT_addr = wIdx[15:0];
  assign MEM_0_MPORT_mask = io_in_wstrb[0];
  assign MEM_0_MPORT_en = _T_42 & _T_52;
  assign MEM_1_MPORT_1_en = 1'h1;
  assign MEM_1_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_1_MPORT_1_data = MEM_1[MEM_1_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_1_MPORT_1_data = MEM_1_MPORT_1_addr >= 16'hea60 ? _RAND_3[7:0] : MEM_1[MEM_1_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_1_MPORT_data = io_in_wdata[15:8];
  assign MEM_1_MPORT_addr = wIdx[15:0];
  assign MEM_1_MPORT_mask = io_in_wstrb[1];
  assign MEM_1_MPORT_en = _T_42 & _T_52;
  assign MEM_2_MPORT_1_en = 1'h1;
  assign MEM_2_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_2_MPORT_1_data = MEM_2[MEM_2_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_2_MPORT_1_data = MEM_2_MPORT_1_addr >= 16'hea60 ? _RAND_5[7:0] : MEM_2[MEM_2_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_2_MPORT_data = io_in_wdata[23:16];
  assign MEM_2_MPORT_addr = wIdx[15:0];
  assign MEM_2_MPORT_mask = io_in_wstrb[2];
  assign MEM_2_MPORT_en = _T_42 & _T_52;
  assign MEM_3_MPORT_1_en = 1'h1;
  assign MEM_3_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_3_MPORT_1_data = MEM_3[MEM_3_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_3_MPORT_1_data = MEM_3_MPORT_1_addr >= 16'hea60 ? _RAND_7[7:0] : MEM_3[MEM_3_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_3_MPORT_data = io_in_wdata[31:24];
  assign MEM_3_MPORT_addr = wIdx[15:0];
  assign MEM_3_MPORT_mask = io_in_wstrb[3];
  assign MEM_3_MPORT_en = _T_42 & _T_52;
  assign MEM_4_MPORT_1_en = 1'h1;
  assign MEM_4_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_4_MPORT_1_data = MEM_4[MEM_4_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_4_MPORT_1_data = MEM_4_MPORT_1_addr >= 16'hea60 ? _RAND_9[7:0] : MEM_4[MEM_4_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_4_MPORT_data = io_in_wdata[39:32];
  assign MEM_4_MPORT_addr = wIdx[15:0];
  assign MEM_4_MPORT_mask = io_in_wstrb[4];
  assign MEM_4_MPORT_en = _T_42 & _T_52;
  assign MEM_5_MPORT_1_en = 1'h1;
  assign MEM_5_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_5_MPORT_1_data = MEM_5[MEM_5_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_5_MPORT_1_data = MEM_5_MPORT_1_addr >= 16'hea60 ? _RAND_11[7:0] : MEM_5[MEM_5_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_5_MPORT_data = io_in_wdata[47:40];
  assign MEM_5_MPORT_addr = wIdx[15:0];
  assign MEM_5_MPORT_mask = io_in_wstrb[5];
  assign MEM_5_MPORT_en = _T_42 & _T_52;
  assign MEM_6_MPORT_1_en = 1'h1;
  assign MEM_6_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_6_MPORT_1_data = MEM_6[MEM_6_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_6_MPORT_1_data = MEM_6_MPORT_1_addr >= 16'hea60 ? _RAND_13[7:0] : MEM_6[MEM_6_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_6_MPORT_data = io_in_wdata[55:48];
  assign MEM_6_MPORT_addr = wIdx[15:0];
  assign MEM_6_MPORT_mask = io_in_wstrb[6];
  assign MEM_6_MPORT_en = _T_42 & _T_52;
  assign MEM_7_MPORT_1_en = 1'h1;
  assign MEM_7_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_7_MPORT_1_data = MEM_7[MEM_7_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_7_MPORT_1_data = MEM_7_MPORT_1_addr >= 16'hea60 ? _RAND_15[7:0] : MEM_7[MEM_7_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_7_MPORT_data = io_in_wdata[63:56];
  assign MEM_7_MPORT_addr = wIdx[15:0];
  assign MEM_7_MPORT_mask = io_in_wstrb[7];
  assign MEM_7_MPORT_en = _T_42 & _T_52;
  assign io_in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io_in_wready = io_in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io_in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io_in_arready = 1'h1; // @[AXI4Slave.scala 71:29]
  assign io_in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io_in_rdata = r; // @[AXI4RAM.scala 71:18]
  always @(posedge clock) begin
    if (MEM_0_MPORT_en & MEM_0_MPORT_mask) begin
      MEM_0[MEM_0_MPORT_addr] <= MEM_0_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_1_MPORT_en & MEM_1_MPORT_mask) begin
      MEM_1[MEM_1_MPORT_addr] <= MEM_1_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_2_MPORT_en & MEM_2_MPORT_mask) begin
      MEM_2[MEM_2_MPORT_addr] <= MEM_2_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_3_MPORT_en & MEM_3_MPORT_mask) begin
      MEM_3[MEM_3_MPORT_addr] <= MEM_3_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_4_MPORT_en & MEM_4_MPORT_mask) begin
      MEM_4[MEM_4_MPORT_addr] <= MEM_4_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_5_MPORT_en & MEM_5_MPORT_mask) begin
      MEM_5[MEM_5_MPORT_addr] <= MEM_5_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_6_MPORT_en & MEM_6_MPORT_mask) begin
      MEM_6[MEM_6_MPORT_addr] <= MEM_6_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_7_MPORT_en & MEM_7_MPORT_mask) begin
      MEM_7[MEM_7_MPORT_addr] <= MEM_7_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    if (REG) begin // @[Reg.scala 16:19]
      r <= rdata; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG_2 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  r = _RAND_21[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_awready,
  input         io_in_fb_awvalid,
  input  [31:0] io_in_fb_awaddr,
  input  [2:0]  io_in_fb_awprot,
  output        io_in_fb_wready,
  input         io_in_fb_wvalid,
  input  [63:0] io_in_fb_wdata,
  input  [7:0]  io_in_fb_wstrb,
  input         io_in_fb_bready,
  output        io_in_fb_bvalid,
  output [1:0]  io_in_fb_bresp,
  output        io_in_fb_arready,
  input         io_in_fb_arvalid,
  input  [31:0] io_in_fb_araddr,
  input  [2:0]  io_in_fb_arprot,
  input         io_in_fb_rready,
  output        io_in_fb_rvalid,
  output [1:0]  io_in_fb_rresp,
  output [63:0] io_in_fb_rdata,
  output        io_in_ctrl_awready,
  input         io_in_ctrl_awvalid,
  input  [31:0] io_in_ctrl_awaddr,
  input  [2:0]  io_in_ctrl_awprot,
  output        io_in_ctrl_wready,
  input         io_in_ctrl_wvalid,
  input  [63:0] io_in_ctrl_wdata,
  input  [7:0]  io_in_ctrl_wstrb,
  input         io_in_ctrl_bready,
  output        io_in_ctrl_bvalid,
  output [1:0]  io_in_ctrl_bresp,
  output        io_in_ctrl_arready,
  input         io_in_ctrl_arvalid,
  input  [31:0] io_in_ctrl_araddr,
  input  [2:0]  io_in_ctrl_arprot,
  input         io_in_ctrl_rready,
  output        io_in_ctrl_rvalid,
  output [1:0]  io_in_ctrl_rresp,
  output [63:0] io_in_ctrl_rdata,
  output [23:0] io_vga_rgb,
  output        io_vga_hsync,
  output        io_vga_vsync,
  output        io_vga_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_awready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_awvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_wready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_wvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_bready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_bvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_arready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_arvalid; // @[AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_araddr; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_rready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_rvalid; // @[AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_rdata; // @[AXI4VGA.scala 125:20]
  wire  fb_clock; // @[AXI4VGA.scala 127:18]
  wire  fb_reset; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_awready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_awvalid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_awaddr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_wready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_wvalid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_wdata; // @[AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_wstrb; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_bready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_bvalid; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_arready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_arvalid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_araddr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_rready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_rvalid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_rdata; // @[AXI4VGA.scala 127:18]
  wire  _T = io_in_fb_arready & io_in_fb_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_1 = io_in_fb_rready & io_in_fb_rvalid; // @[Decoupled.scala 40:37]
  reg  REG; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_1 ? 1'h0 : REG; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg [10:0] hCounter; // @[Counter.scala 60:40]
  wire  wrap_wrap = hCounter == 11'h41f; // @[Counter.scala 72:24]
  wire [10:0] _wrap_value_T_1 = hCounter + 11'h1; // @[Counter.scala 76:24]
  reg [9:0] vCounter; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = vCounter == 10'h273; // @[Counter.scala 72:24]
  wire [9:0] _wrap_value_T_3 = vCounter + 10'h1; // @[Counter.scala 76:24]
  wire  hInRange = hCounter >= 11'ha8 & hCounter < 11'h3c8; // @[AXI4VGA.scala 138:63]
  wire  vInRange = vCounter >= 10'h5 & vCounter < 10'h25d; // @[AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[AXI4VGA.scala 152:31]
  wire  _T_12 = hCounter >= 11'ha7 & hCounter < 11'h3c7; // @[AXI4VGA.scala 138:63]
  wire  nextPixel = _T_12 & vInRange & hCounterIsOdd; // @[AXI4VGA.scala 155:78]
  wire  _T_15 = nextPixel & ~vCounterIsOdd; // @[AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[Counter.scala 60:40]
  wire  wrap_wrap_2 = fbPixelAddrV0 == 17'h1d4bf; // @[Counter.scala 72:24]
  wire [16:0] _wrap_value_T_5 = fbPixelAddrV0 + 17'h1; // @[Counter.scala 76:24]
  wire  _T_16 = nextPixel & vCounterIsOdd; // @[AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[Counter.scala 60:40]
  wire  wrap_wrap_3 = fbPixelAddrV1 == 17'h1d4bf; // @[Counter.scala 72:24]
  wire [16:0] _wrap_value_T_7 = fbPixelAddrV1 + 17'h1; // @[Counter.scala 76:24]
  wire [16:0] _T_17 = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[AXI4VGA.scala 161:35]
  wire [18:0] _T_18 = {_T_17,2'h0}; // @[Cat.scala 30:58]
  reg  REG_1; // @[AXI4VGA.scala 162:31]
  wire  _T_20 = fb_io_in_rready & fb_io_in_rvalid; // @[Decoupled.scala 40:37]
  reg [63:0] r; // @[Reg.scala 27:20]
  wire [63:0] _GEN_14 = _T_20 ? fb_io_in_rdata : r; // @[Reg.scala 28:19 27:20 28:23]
  wire [31:0] color = hCounter[1] ? _GEN_14[63:32] : _GEN_14[31:0]; // @[AXI4VGA.scala 167:23]
  VGACtrl ctrl ( // @[AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_awready(ctrl_io_in_awready),
    .io_in_awvalid(ctrl_io_in_awvalid),
    .io_in_wready(ctrl_io_in_wready),
    .io_in_wvalid(ctrl_io_in_wvalid),
    .io_in_bready(ctrl_io_in_bready),
    .io_in_bvalid(ctrl_io_in_bvalid),
    .io_in_arready(ctrl_io_in_arready),
    .io_in_arvalid(ctrl_io_in_arvalid),
    .io_in_araddr(ctrl_io_in_araddr),
    .io_in_rready(ctrl_io_in_rready),
    .io_in_rvalid(ctrl_io_in_rvalid),
    .io_in_rdata(ctrl_io_in_rdata)
  );
  AXI4RAM fb ( // @[AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_awready(fb_io_in_awready),
    .io_in_awvalid(fb_io_in_awvalid),
    .io_in_awaddr(fb_io_in_awaddr),
    .io_in_wready(fb_io_in_wready),
    .io_in_wvalid(fb_io_in_wvalid),
    .io_in_wdata(fb_io_in_wdata),
    .io_in_wstrb(fb_io_in_wstrb),
    .io_in_bready(fb_io_in_bready),
    .io_in_bvalid(fb_io_in_bvalid),
    .io_in_arready(fb_io_in_arready),
    .io_in_arvalid(fb_io_in_arvalid),
    .io_in_araddr(fb_io_in_araddr),
    .io_in_rready(fb_io_in_rready),
    .io_in_rvalid(fb_io_in_rvalid),
    .io_in_rdata(fb_io_in_rdata)
  );
  assign io_in_fb_awready = fb_io_in_awready; // @[AXI4VGA.scala 130:15]
  assign io_in_fb_wready = fb_io_in_wready; // @[AXI4VGA.scala 131:14]
  assign io_in_fb_bvalid = fb_io_in_bvalid; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_bresp = 2'h0; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_arready = 1'h1; // @[AXI4VGA.scala 133:21]
  assign io_in_fb_rvalid = REG; // @[AXI4VGA.scala 136:20]
  assign io_in_fb_rresp = 2'h0; // @[AXI4VGA.scala 135:24]
  assign io_in_fb_rdata = 64'h0; // @[AXI4VGA.scala 134:24]
  assign io_in_ctrl_awready = ctrl_io_in_awready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_wready = ctrl_io_in_wready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_bvalid = ctrl_io_in_bvalid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_bresp = 2'h0; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_arready = ctrl_io_in_arready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rvalid = ctrl_io_in_rvalid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rresp = 2'h0; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rdata = ctrl_io_in_rdata; // @[AXI4VGA.scala 126:14]
  assign io_vga_rgb = io_vga_valid ? color[23:0] : 24'h0; // @[AXI4VGA.scala 168:20]
  assign io_vga_hsync = hCounter >= 11'h28; // @[AXI4VGA.scala 143:28]
  assign io_vga_vsync = vCounter >= 10'h1; // @[AXI4VGA.scala 144:28]
  assign io_vga_valid = hInRange & vInRange; // @[AXI4VGA.scala 148:28]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_awvalid = io_in_ctrl_awvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_wvalid = io_in_ctrl_wvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_bready = io_in_ctrl_bready; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_arvalid = io_in_ctrl_arvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_araddr = io_in_ctrl_araddr; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_rready = io_in_ctrl_rready; // @[AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_awvalid = io_in_fb_awvalid; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_awaddr = io_in_fb_awaddr; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_wvalid = io_in_fb_wvalid; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_wdata = io_in_fb_wdata; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_wstrb = io_in_fb_wstrb; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_bready = io_in_fb_bready; // @[AXI4VGA.scala 132:14]
  assign fb_io_in_arvalid = REG_1 & hCounterIs2; // @[AXI4VGA.scala 162:43]
  assign fb_io_in_araddr = {{13'd0}, _T_18}; // @[AXI4VGA.scala 161:25]
  assign fb_io_in_rready = 1'h1; // @[AXI4VGA.scala 164:20]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      REG <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG <= _GEN_1;
    end
    if (reset) begin // @[Counter.scala 60:40]
      hCounter <= 11'h0; // @[Counter.scala 60:40]
    end else if (wrap_wrap) begin // @[Counter.scala 86:20]
      hCounter <= 11'h0; // @[Counter.scala 86:28]
    end else begin
      hCounter <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      vCounter <= 10'h0; // @[Counter.scala 60:40]
    end else if (wrap_wrap) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        vCounter <= 10'h0; // @[Counter.scala 86:28]
      end else begin
        vCounter <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      fbPixelAddrV0 <= 17'h0; // @[Counter.scala 60:40]
    end else if (_T_15) begin // @[Counter.scala 118:17]
      if (wrap_wrap_2) begin // @[Counter.scala 86:20]
        fbPixelAddrV0 <= 17'h0; // @[Counter.scala 86:28]
      end else begin
        fbPixelAddrV0 <= _wrap_value_T_5; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      fbPixelAddrV1 <= 17'h0; // @[Counter.scala 60:40]
    end else if (_T_16) begin // @[Counter.scala 118:17]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20]
        fbPixelAddrV1 <= 17'h0; // @[Counter.scala 86:28]
      end else begin
        fbPixelAddrV1 <= _wrap_value_T_7; // @[Counter.scala 76:15]
      end
    end
    REG_1 <= _T_12 & vInRange & hCounterIsOdd; // @[AXI4VGA.scala 155:78]
    if (reset) begin // @[Reg.scala 27:20]
      r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      r <= fb_io_in_rdata; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hCounter = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  vCounter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input   clock,
  input   reset
);
  wire  nutshell_clock; // @[TopMain.scala 29:24]
  wire  nutshell_reset; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mem_awaddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_awprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awuser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mem_awlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_awsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_awburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_awcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_awqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_wready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_wvalid; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mem_wdata; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mem_wstrb; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_wlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_bready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_bvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_bresp; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_bid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_buser; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mem_araddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_arprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_aruser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mem_arlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_arsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_arburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_arcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_arqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_rresp; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mem_rdata; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_ruser; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mmio_awaddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_awprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awuser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mmio_awlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_awsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_awburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_awcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_awqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_wready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_wvalid; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mmio_wdata; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mmio_wstrb; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_wlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_bready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_bvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_bresp; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_bid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_buser; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mmio_araddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_arprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_aruser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mmio_arlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_arsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_arburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_arcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_arqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_rresp; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mmio_rdata; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_ruser; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_frontend_awaddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_awprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awuser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_frontend_awlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_awsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_awburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_awcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_awqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_wready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_wvalid; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_frontend_wdata; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_frontend_wstrb; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_wlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_bready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_bvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_bresp; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_bid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_buser; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_frontend_araddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_arprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_aruser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_frontend_arlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_arsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_arburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_arcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_arqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_rresp; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_frontend_rdata; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_ruser; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_meip; // @[TopMain.scala 29:24]
  wire [38:0] nutshell_io_ila_WBUpc; // @[TopMain.scala 29:24]
  wire  nutshell_io_ila_WBUvalid; // @[TopMain.scala 29:24]
  wire  nutshell_io_ila_WBUrfWen; // @[TopMain.scala 29:24]
  wire [4:0] nutshell_io_ila_WBUrfDest; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_ila_WBUrfData; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_ila_InstrCnt; // @[TopMain.scala 29:24]
  wire  vga_clock; // @[TopMain.scala 30:19]
  wire  vga_reset; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_awready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_awvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_fb_awaddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_fb_awprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_wready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_wvalid; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_fb_wdata; // @[TopMain.scala 30:19]
  wire [7:0] vga_io_in_fb_wstrb; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_bready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_bvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_fb_bresp; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_arready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_arvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_fb_araddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_fb_arprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_rready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_rvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_fb_rresp; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_fb_rdata; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_awready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_awvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_ctrl_awaddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_ctrl_awprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_wready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_wvalid; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_ctrl_wdata; // @[TopMain.scala 30:19]
  wire [7:0] vga_io_in_ctrl_wstrb; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_bready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_bvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_ctrl_bresp; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_arready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_arvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_ctrl_araddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_ctrl_arprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_rready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_rvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_ctrl_rresp; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_ctrl_rdata; // @[TopMain.scala 30:19]
  wire [23:0] vga_io_vga_rgb; // @[TopMain.scala 30:19]
  wire  vga_io_vga_hsync; // @[TopMain.scala 30:19]
  wire  vga_io_vga_vsync; // @[TopMain.scala 30:19]
  wire  vga_io_vga_valid; // @[TopMain.scala 30:19]
  NutShell nutshell ( // @[TopMain.scala 29:24]
    .clock(nutshell_clock),
    .reset(nutshell_reset),
    .io_mem_awready(nutshell_io_mem_awready),
    .io_mem_awvalid(nutshell_io_mem_awvalid),
    .io_mem_awaddr(nutshell_io_mem_awaddr),
    .io_mem_awprot(nutshell_io_mem_awprot),
    .io_mem_awid(nutshell_io_mem_awid),
    .io_mem_awuser(nutshell_io_mem_awuser),
    .io_mem_awlen(nutshell_io_mem_awlen),
    .io_mem_awsize(nutshell_io_mem_awsize),
    .io_mem_awburst(nutshell_io_mem_awburst),
    .io_mem_awlock(nutshell_io_mem_awlock),
    .io_mem_awcache(nutshell_io_mem_awcache),
    .io_mem_awqos(nutshell_io_mem_awqos),
    .io_mem_wready(nutshell_io_mem_wready),
    .io_mem_wvalid(nutshell_io_mem_wvalid),
    .io_mem_wdata(nutshell_io_mem_wdata),
    .io_mem_wstrb(nutshell_io_mem_wstrb),
    .io_mem_wlast(nutshell_io_mem_wlast),
    .io_mem_bready(nutshell_io_mem_bready),
    .io_mem_bvalid(nutshell_io_mem_bvalid),
    .io_mem_bresp(nutshell_io_mem_bresp),
    .io_mem_bid(nutshell_io_mem_bid),
    .io_mem_buser(nutshell_io_mem_buser),
    .io_mem_arready(nutshell_io_mem_arready),
    .io_mem_arvalid(nutshell_io_mem_arvalid),
    .io_mem_araddr(nutshell_io_mem_araddr),
    .io_mem_arprot(nutshell_io_mem_arprot),
    .io_mem_arid(nutshell_io_mem_arid),
    .io_mem_aruser(nutshell_io_mem_aruser),
    .io_mem_arlen(nutshell_io_mem_arlen),
    .io_mem_arsize(nutshell_io_mem_arsize),
    .io_mem_arburst(nutshell_io_mem_arburst),
    .io_mem_arlock(nutshell_io_mem_arlock),
    .io_mem_arcache(nutshell_io_mem_arcache),
    .io_mem_arqos(nutshell_io_mem_arqos),
    .io_mem_rready(nutshell_io_mem_rready),
    .io_mem_rvalid(nutshell_io_mem_rvalid),
    .io_mem_rresp(nutshell_io_mem_rresp),
    .io_mem_rdata(nutshell_io_mem_rdata),
    .io_mem_rlast(nutshell_io_mem_rlast),
    .io_mem_rid(nutshell_io_mem_rid),
    .io_mem_ruser(nutshell_io_mem_ruser),
    .io_mmio_awready(nutshell_io_mmio_awready),
    .io_mmio_awvalid(nutshell_io_mmio_awvalid),
    .io_mmio_awaddr(nutshell_io_mmio_awaddr),
    .io_mmio_awprot(nutshell_io_mmio_awprot),
    .io_mmio_awid(nutshell_io_mmio_awid),
    .io_mmio_awuser(nutshell_io_mmio_awuser),
    .io_mmio_awlen(nutshell_io_mmio_awlen),
    .io_mmio_awsize(nutshell_io_mmio_awsize),
    .io_mmio_awburst(nutshell_io_mmio_awburst),
    .io_mmio_awlock(nutshell_io_mmio_awlock),
    .io_mmio_awcache(nutshell_io_mmio_awcache),
    .io_mmio_awqos(nutshell_io_mmio_awqos),
    .io_mmio_wready(nutshell_io_mmio_wready),
    .io_mmio_wvalid(nutshell_io_mmio_wvalid),
    .io_mmio_wdata(nutshell_io_mmio_wdata),
    .io_mmio_wstrb(nutshell_io_mmio_wstrb),
    .io_mmio_wlast(nutshell_io_mmio_wlast),
    .io_mmio_bready(nutshell_io_mmio_bready),
    .io_mmio_bvalid(nutshell_io_mmio_bvalid),
    .io_mmio_bresp(nutshell_io_mmio_bresp),
    .io_mmio_bid(nutshell_io_mmio_bid),
    .io_mmio_buser(nutshell_io_mmio_buser),
    .io_mmio_arready(nutshell_io_mmio_arready),
    .io_mmio_arvalid(nutshell_io_mmio_arvalid),
    .io_mmio_araddr(nutshell_io_mmio_araddr),
    .io_mmio_arprot(nutshell_io_mmio_arprot),
    .io_mmio_arid(nutshell_io_mmio_arid),
    .io_mmio_aruser(nutshell_io_mmio_aruser),
    .io_mmio_arlen(nutshell_io_mmio_arlen),
    .io_mmio_arsize(nutshell_io_mmio_arsize),
    .io_mmio_arburst(nutshell_io_mmio_arburst),
    .io_mmio_arlock(nutshell_io_mmio_arlock),
    .io_mmio_arcache(nutshell_io_mmio_arcache),
    .io_mmio_arqos(nutshell_io_mmio_arqos),
    .io_mmio_rready(nutshell_io_mmio_rready),
    .io_mmio_rvalid(nutshell_io_mmio_rvalid),
    .io_mmio_rresp(nutshell_io_mmio_rresp),
    .io_mmio_rdata(nutshell_io_mmio_rdata),
    .io_mmio_rlast(nutshell_io_mmio_rlast),
    .io_mmio_rid(nutshell_io_mmio_rid),
    .io_mmio_ruser(nutshell_io_mmio_ruser),
    .io_frontend_awready(nutshell_io_frontend_awready),
    .io_frontend_awvalid(nutshell_io_frontend_awvalid),
    .io_frontend_awaddr(nutshell_io_frontend_awaddr),
    .io_frontend_awprot(nutshell_io_frontend_awprot),
    .io_frontend_awid(nutshell_io_frontend_awid),
    .io_frontend_awuser(nutshell_io_frontend_awuser),
    .io_frontend_awlen(nutshell_io_frontend_awlen),
    .io_frontend_awsize(nutshell_io_frontend_awsize),
    .io_frontend_awburst(nutshell_io_frontend_awburst),
    .io_frontend_awlock(nutshell_io_frontend_awlock),
    .io_frontend_awcache(nutshell_io_frontend_awcache),
    .io_frontend_awqos(nutshell_io_frontend_awqos),
    .io_frontend_wready(nutshell_io_frontend_wready),
    .io_frontend_wvalid(nutshell_io_frontend_wvalid),
    .io_frontend_wdata(nutshell_io_frontend_wdata),
    .io_frontend_wstrb(nutshell_io_frontend_wstrb),
    .io_frontend_wlast(nutshell_io_frontend_wlast),
    .io_frontend_bready(nutshell_io_frontend_bready),
    .io_frontend_bvalid(nutshell_io_frontend_bvalid),
    .io_frontend_bresp(nutshell_io_frontend_bresp),
    .io_frontend_bid(nutshell_io_frontend_bid),
    .io_frontend_buser(nutshell_io_frontend_buser),
    .io_frontend_arready(nutshell_io_frontend_arready),
    .io_frontend_arvalid(nutshell_io_frontend_arvalid),
    .io_frontend_araddr(nutshell_io_frontend_araddr),
    .io_frontend_arprot(nutshell_io_frontend_arprot),
    .io_frontend_arid(nutshell_io_frontend_arid),
    .io_frontend_aruser(nutshell_io_frontend_aruser),
    .io_frontend_arlen(nutshell_io_frontend_arlen),
    .io_frontend_arsize(nutshell_io_frontend_arsize),
    .io_frontend_arburst(nutshell_io_frontend_arburst),
    .io_frontend_arlock(nutshell_io_frontend_arlock),
    .io_frontend_arcache(nutshell_io_frontend_arcache),
    .io_frontend_arqos(nutshell_io_frontend_arqos),
    .io_frontend_rready(nutshell_io_frontend_rready),
    .io_frontend_rvalid(nutshell_io_frontend_rvalid),
    .io_frontend_rresp(nutshell_io_frontend_rresp),
    .io_frontend_rdata(nutshell_io_frontend_rdata),
    .io_frontend_rlast(nutshell_io_frontend_rlast),
    .io_frontend_rid(nutshell_io_frontend_rid),
    .io_frontend_ruser(nutshell_io_frontend_ruser),
    .io_meip(nutshell_io_meip),
    .io_ila_WBUpc(nutshell_io_ila_WBUpc),
    .io_ila_WBUvalid(nutshell_io_ila_WBUvalid),
    .io_ila_WBUrfWen(nutshell_io_ila_WBUrfWen),
    .io_ila_WBUrfDest(nutshell_io_ila_WBUrfDest),
    .io_ila_WBUrfData(nutshell_io_ila_WBUrfData),
    .io_ila_InstrCnt(nutshell_io_ila_InstrCnt)
  );
  AXI4VGA vga ( // @[TopMain.scala 30:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_awready(vga_io_in_fb_awready),
    .io_in_fb_awvalid(vga_io_in_fb_awvalid),
    .io_in_fb_awaddr(vga_io_in_fb_awaddr),
    .io_in_fb_awprot(vga_io_in_fb_awprot),
    .io_in_fb_wready(vga_io_in_fb_wready),
    .io_in_fb_wvalid(vga_io_in_fb_wvalid),
    .io_in_fb_wdata(vga_io_in_fb_wdata),
    .io_in_fb_wstrb(vga_io_in_fb_wstrb),
    .io_in_fb_bready(vga_io_in_fb_bready),
    .io_in_fb_bvalid(vga_io_in_fb_bvalid),
    .io_in_fb_bresp(vga_io_in_fb_bresp),
    .io_in_fb_arready(vga_io_in_fb_arready),
    .io_in_fb_arvalid(vga_io_in_fb_arvalid),
    .io_in_fb_araddr(vga_io_in_fb_araddr),
    .io_in_fb_arprot(vga_io_in_fb_arprot),
    .io_in_fb_rready(vga_io_in_fb_rready),
    .io_in_fb_rvalid(vga_io_in_fb_rvalid),
    .io_in_fb_rresp(vga_io_in_fb_rresp),
    .io_in_fb_rdata(vga_io_in_fb_rdata),
    .io_in_ctrl_awready(vga_io_in_ctrl_awready),
    .io_in_ctrl_awvalid(vga_io_in_ctrl_awvalid),
    .io_in_ctrl_awaddr(vga_io_in_ctrl_awaddr),
    .io_in_ctrl_awprot(vga_io_in_ctrl_awprot),
    .io_in_ctrl_wready(vga_io_in_ctrl_wready),
    .io_in_ctrl_wvalid(vga_io_in_ctrl_wvalid),
    .io_in_ctrl_wdata(vga_io_in_ctrl_wdata),
    .io_in_ctrl_wstrb(vga_io_in_ctrl_wstrb),
    .io_in_ctrl_bready(vga_io_in_ctrl_bready),
    .io_in_ctrl_bvalid(vga_io_in_ctrl_bvalid),
    .io_in_ctrl_bresp(vga_io_in_ctrl_bresp),
    .io_in_ctrl_arready(vga_io_in_ctrl_arready),
    .io_in_ctrl_arvalid(vga_io_in_ctrl_arvalid),
    .io_in_ctrl_araddr(vga_io_in_ctrl_araddr),
    .io_in_ctrl_arprot(vga_io_in_ctrl_arprot),
    .io_in_ctrl_rready(vga_io_in_ctrl_rready),
    .io_in_ctrl_rvalid(vga_io_in_ctrl_rvalid),
    .io_in_ctrl_rresp(vga_io_in_ctrl_rresp),
    .io_in_ctrl_rdata(vga_io_in_ctrl_rdata),
    .io_vga_rgb(vga_io_vga_rgb),
    .io_vga_hsync(vga_io_vga_hsync),
    .io_vga_vsync(vga_io_vga_vsync),
    .io_vga_valid(vga_io_vga_valid)
  );
  assign nutshell_clock = clock;
  assign nutshell_reset = reset;
  assign nutshell_io_mem_awready = 1'h0;
  assign nutshell_io_mem_wready = 1'h0;
  assign nutshell_io_mem_bvalid = 1'h0;
  assign nutshell_io_mem_bresp = 2'h0;
  assign nutshell_io_mem_bid = 1'h0;
  assign nutshell_io_mem_buser = 1'h0;
  assign nutshell_io_mem_arready = 1'h0;
  assign nutshell_io_mem_rvalid = 1'h0;
  assign nutshell_io_mem_rresp = 2'h0;
  assign nutshell_io_mem_rdata = 64'h0;
  assign nutshell_io_mem_rlast = 1'h0;
  assign nutshell_io_mem_rid = 1'h0;
  assign nutshell_io_mem_ruser = 1'h0;
  assign nutshell_io_mmio_awready = 1'h0;
  assign nutshell_io_mmio_wready = 1'h0;
  assign nutshell_io_mmio_bvalid = 1'h0;
  assign nutshell_io_mmio_bresp = 2'h0;
  assign nutshell_io_mmio_bid = 1'h0;
  assign nutshell_io_mmio_buser = 1'h0;
  assign nutshell_io_mmio_arready = 1'h0;
  assign nutshell_io_mmio_rvalid = 1'h0;
  assign nutshell_io_mmio_rresp = 2'h0;
  assign nutshell_io_mmio_rdata = 64'h0;
  assign nutshell_io_mmio_rlast = 1'h0;
  assign nutshell_io_mmio_rid = 1'h0;
  assign nutshell_io_mmio_ruser = 1'h0;
  assign nutshell_io_frontend_awvalid = 1'h0;
  assign nutshell_io_frontend_awaddr = 32'h0;
  assign nutshell_io_frontend_awprot = 3'h0;
  assign nutshell_io_frontend_awid = 1'h0;
  assign nutshell_io_frontend_awuser = 1'h0;
  assign nutshell_io_frontend_awlen = 8'h0;
  assign nutshell_io_frontend_awsize = 3'h0;
  assign nutshell_io_frontend_awburst = 2'h0;
  assign nutshell_io_frontend_awlock = 1'h0;
  assign nutshell_io_frontend_awcache = 4'h0;
  assign nutshell_io_frontend_awqos = 4'h0;
  assign nutshell_io_frontend_wvalid = 1'h0;
  assign nutshell_io_frontend_wdata = 64'h0;
  assign nutshell_io_frontend_wstrb = 8'h0;
  assign nutshell_io_frontend_wlast = 1'h0;
  assign nutshell_io_frontend_bready = 1'h0;
  assign nutshell_io_frontend_arvalid = 1'h0;
  assign nutshell_io_frontend_araddr = 32'h0;
  assign nutshell_io_frontend_arprot = 3'h0;
  assign nutshell_io_frontend_arid = 1'h0;
  assign nutshell_io_frontend_aruser = 1'h0;
  assign nutshell_io_frontend_arlen = 8'h0;
  assign nutshell_io_frontend_arsize = 3'h0;
  assign nutshell_io_frontend_arburst = 2'h0;
  assign nutshell_io_frontend_arlock = 1'h0;
  assign nutshell_io_frontend_arcache = 4'h0;
  assign nutshell_io_frontend_arqos = 4'h0;
  assign nutshell_io_frontend_rready = 1'h0;
  assign nutshell_io_meip = 3'h0;
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_awvalid = 1'h0;
  assign vga_io_in_fb_awaddr = 32'h0;
  assign vga_io_in_fb_awprot = 3'h0;
  assign vga_io_in_fb_wvalid = 1'h0;
  assign vga_io_in_fb_wdata = 64'h0;
  assign vga_io_in_fb_wstrb = 8'h0;
  assign vga_io_in_fb_bready = 1'h0;
  assign vga_io_in_fb_arvalid = 1'h0;
  assign vga_io_in_fb_araddr = 32'h0;
  assign vga_io_in_fb_arprot = 3'h0;
  assign vga_io_in_fb_rready = 1'h0;
  assign vga_io_in_ctrl_awvalid = 1'h0;
  assign vga_io_in_ctrl_awaddr = 32'h0;
  assign vga_io_in_ctrl_awprot = 3'h0;
  assign vga_io_in_ctrl_wvalid = 1'h0;
  assign vga_io_in_ctrl_wdata = 64'h0;
  assign vga_io_in_ctrl_wstrb = 8'h0;
  assign vga_io_in_ctrl_bready = 1'h0;
  assign vga_io_in_ctrl_arvalid = 1'h0;
  assign vga_io_in_ctrl_araddr = 32'h0;
  assign vga_io_in_ctrl_arprot = 3'h0;
  assign vga_io_in_ctrl_rready = 1'h0;
endmodule
module array(
  input  [8:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [72:0] RW0_wdata_0,
  output [72:0] RW0_rdata_0
);
  wire [8:0] array_ext_RW0_addr;
  wire  array_ext_RW0_en;
  wire  array_ext_RW0_clk;
  wire  array_ext_RW0_wmode;
  wire [72:0] array_ext_RW0_wdata;
  wire [72:0] array_ext_RW0_rdata;
  array_ext array_ext (
    .RW0_addr(array_ext_RW0_addr),
    .RW0_en(array_ext_RW0_en),
    .RW0_clk(array_ext_RW0_clk),
    .RW0_wmode(array_ext_RW0_wmode),
    .RW0_wdata(array_ext_RW0_wdata),
    .RW0_rdata(array_ext_RW0_rdata)
  );
  assign array_ext_RW0_clk = RW0_clk;
  assign array_ext_RW0_en = RW0_en;
  assign array_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_ext_RW0_rdata;
  assign array_ext_RW0_wmode = RW0_wmode;
  assign array_ext_RW0_wdata = RW0_wdata_0;
endmodule
module array_0(
  input  [6:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [20:0] RW0_wdata_0,
  input  [20:0] RW0_wdata_1,
  input  [20:0] RW0_wdata_2,
  input  [20:0] RW0_wdata_3,
  output [20:0] RW0_rdata_0,
  output [20:0] RW0_rdata_1,
  output [20:0] RW0_rdata_2,
  output [20:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [6:0] array_0_ext_RW0_addr;
  wire  array_0_ext_RW0_en;
  wire  array_0_ext_RW0_clk;
  wire  array_0_ext_RW0_wmode;
  wire [83:0] array_0_ext_RW0_wdata;
  wire [83:0] array_0_ext_RW0_rdata;
  wire [3:0] array_0_ext_RW0_wmask;
  wire [41:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [41:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_0_ext array_0_ext (
    .RW0_addr(array_0_ext_RW0_addr),
    .RW0_en(array_0_ext_RW0_en),
    .RW0_clk(array_0_ext_RW0_clk),
    .RW0_wmode(array_0_ext_RW0_wmode),
    .RW0_wdata(array_0_ext_RW0_wdata),
    .RW0_rdata(array_0_ext_RW0_rdata),
    .RW0_wmask(array_0_ext_RW0_wmask)
  );
  assign array_0_ext_RW0_clk = RW0_clk;
  assign array_0_ext_RW0_en = RW0_en;
  assign array_0_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_0_ext_RW0_rdata[20:0];
  assign RW0_rdata_1 = array_0_ext_RW0_rdata[41:21];
  assign RW0_rdata_2 = array_0_ext_RW0_rdata[62:42];
  assign RW0_rdata_3 = array_0_ext_RW0_rdata[83:63];
  assign array_0_ext_RW0_wmode = RW0_wmode;
  assign array_0_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_0_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_1(
  input  [9:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [63:0] RW0_wdata_0,
  input  [63:0] RW0_wdata_1,
  input  [63:0] RW0_wdata_2,
  input  [63:0] RW0_wdata_3,
  output [63:0] RW0_rdata_0,
  output [63:0] RW0_rdata_1,
  output [63:0] RW0_rdata_2,
  output [63:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [9:0] array_1_ext_RW0_addr;
  wire  array_1_ext_RW0_en;
  wire  array_1_ext_RW0_clk;
  wire  array_1_ext_RW0_wmode;
  wire [255:0] array_1_ext_RW0_wdata;
  wire [255:0] array_1_ext_RW0_rdata;
  wire [3:0] array_1_ext_RW0_wmask;
  wire [127:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [127:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_1_ext array_1_ext (
    .RW0_addr(array_1_ext_RW0_addr),
    .RW0_en(array_1_ext_RW0_en),
    .RW0_clk(array_1_ext_RW0_clk),
    .RW0_wmode(array_1_ext_RW0_wmode),
    .RW0_wdata(array_1_ext_RW0_wdata),
    .RW0_rdata(array_1_ext_RW0_rdata),
    .RW0_wmask(array_1_ext_RW0_wmask)
  );
  assign array_1_ext_RW0_clk = RW0_clk;
  assign array_1_ext_RW0_en = RW0_en;
  assign array_1_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_1_ext_RW0_rdata[63:0];
  assign RW0_rdata_1 = array_1_ext_RW0_rdata[127:64];
  assign RW0_rdata_2 = array_1_ext_RW0_rdata[191:128];
  assign RW0_rdata_3 = array_1_ext_RW0_rdata[255:192];
  assign array_1_ext_RW0_wmode = RW0_wmode;
  assign array_1_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_1_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_2(
  input  [8:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [18:0] RW0_wdata_0,
  input  [18:0] RW0_wdata_1,
  input  [18:0] RW0_wdata_2,
  input  [18:0] RW0_wdata_3,
  output [18:0] RW0_rdata_0,
  output [18:0] RW0_rdata_1,
  output [18:0] RW0_rdata_2,
  output [18:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [8:0] array_2_ext_RW0_addr;
  wire  array_2_ext_RW0_en;
  wire  array_2_ext_RW0_clk;
  wire  array_2_ext_RW0_wmode;
  wire [75:0] array_2_ext_RW0_wdata;
  wire [75:0] array_2_ext_RW0_rdata;
  wire [3:0] array_2_ext_RW0_wmask;
  wire [37:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [37:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_2_ext array_2_ext (
    .RW0_addr(array_2_ext_RW0_addr),
    .RW0_en(array_2_ext_RW0_en),
    .RW0_clk(array_2_ext_RW0_clk),
    .RW0_wmode(array_2_ext_RW0_wmode),
    .RW0_wdata(array_2_ext_RW0_wdata),
    .RW0_rdata(array_2_ext_RW0_rdata),
    .RW0_wmask(array_2_ext_RW0_wmask)
  );
  assign array_2_ext_RW0_clk = RW0_clk;
  assign array_2_ext_RW0_en = RW0_en;
  assign array_2_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_2_ext_RW0_rdata[18:0];
  assign RW0_rdata_1 = array_2_ext_RW0_rdata[37:19];
  assign RW0_rdata_2 = array_2_ext_RW0_rdata[56:38];
  assign RW0_rdata_3 = array_2_ext_RW0_rdata[75:57];
  assign array_2_ext_RW0_wmode = RW0_wmode;
  assign array_2_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_2_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_3(
  input  [11:0] RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [63:0] RW0_wdata_0,
  input  [63:0] RW0_wdata_1,
  input  [63:0] RW0_wdata_2,
  input  [63:0] RW0_wdata_3,
  output [63:0] RW0_rdata_0,
  output [63:0] RW0_rdata_1,
  output [63:0] RW0_rdata_2,
  output [63:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [11:0] array_3_ext_RW0_addr;
  wire  array_3_ext_RW0_en;
  wire  array_3_ext_RW0_clk;
  wire  array_3_ext_RW0_wmode;
  wire [255:0] array_3_ext_RW0_wdata;
  wire [255:0] array_3_ext_RW0_rdata;
  wire [3:0] array_3_ext_RW0_wmask;
  wire [127:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [127:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_3_ext array_3_ext (
    .RW0_addr(array_3_ext_RW0_addr),
    .RW0_en(array_3_ext_RW0_en),
    .RW0_clk(array_3_ext_RW0_clk),
    .RW0_wmode(array_3_ext_RW0_wmode),
    .RW0_wdata(array_3_ext_RW0_wdata),
    .RW0_rdata(array_3_ext_RW0_rdata),
    .RW0_wmask(array_3_ext_RW0_wmask)
  );
  assign array_3_ext_RW0_clk = RW0_clk;
  assign array_3_ext_RW0_en = RW0_en;
  assign array_3_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_3_ext_RW0_rdata[63:0];
  assign RW0_rdata_1 = array_3_ext_RW0_rdata[127:64];
  assign RW0_rdata_2 = array_3_ext_RW0_rdata[191:128];
  assign RW0_rdata_3 = array_3_ext_RW0_rdata[255:192];
  assign array_3_ext_RW0_wmode = RW0_wmode;
  assign array_3_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_3_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
